`timescale 1ns / 1ps
`include "macro.vh"
///////////////////////
module FIFO( in , out , clk ,reset);

input  [`DATA_LENGTH-1:0] in;
output [`DATA_LENGTH-1:0] out;
input  clk ,reset;
reg	[`DATA_LENGTH-1:0] fifo [0:`W-1];

assign  out =  fifo[`W-1] ;
always @(posedge clk)
begin
	if(reset)
	begin
		fifo[0] <= 0;
		fifo[1] <= 0;
		fifo[2] <= 0;
		fifo[3] <= 0;
		fifo[4] <= 0;
		fifo[5] <= 0;
		fifo[6] <= 0;
		fifo[7] <= 0;
		fifo[8] <= 0;
		fifo[9] <= 0;
		fifo[10] <= 0;
		fifo[11] <= 0;
		fifo[12] <= 0;
		fifo[13] <= 0;
		fifo[14] <= 0;
		fifo[15] <= 0;
		fifo[16] <= 0;
		fifo[17] <= 0;
		fifo[18] <= 0;
		fifo[19] <= 0;
		fifo[20] <= 0;
		fifo[21] <= 0;
		fifo[22] <= 0;
		fifo[23] <= 0;
		fifo[24] <= 0;
		fifo[25] <= 0;
		fifo[26] <= 0;
		fifo[27] <= 0;
		fifo[28] <= 0;
		fifo[29] <= 0;
		fifo[30] <= 0;
		fifo[31] <= 0;
		fifo[32] <= 0;
		fifo[33] <= 0;
		fifo[34] <= 0;
		fifo[35] <= 0;
		fifo[36] <= 0;
		fifo[37] <= 0;
		fifo[38] <= 0;
		fifo[39] <= 0;
		fifo[40] <= 0;
		fifo[41] <= 0;
		fifo[42] <= 0;
		fifo[43] <= 0;
		fifo[44] <= 0;
		fifo[45] <= 0;
		fifo[46] <= 0;
		fifo[47] <= 0;
		fifo[48] <= 0;
		fifo[49] <= 0;
		fifo[50] <= 0;
		fifo[51] <= 0;
		fifo[52] <= 0;
		fifo[53] <= 0;
		fifo[54] <= 0;
		fifo[55] <= 0;
		fifo[56] <= 0;
		fifo[57] <= 0;
		fifo[58] <= 0;
		fifo[59] <= 0;
		fifo[60] <= 0;
		fifo[61] <= 0;
		fifo[62] <= 0;
		fifo[63] <= 0;
		fifo[64] <= 0;
		fifo[65] <= 0;
		fifo[66] <= 0;
		fifo[67] <= 0;
		fifo[68] <= 0;
		fifo[69] <= 0;
		fifo[70] <= 0;
		fifo[71] <= 0;
		fifo[72] <= 0;
		fifo[73] <= 0;
		fifo[74] <= 0;
		fifo[75] <= 0;
		fifo[76] <= 0;
		fifo[77] <= 0;
		fifo[78] <= 0;
		fifo[79] <= 0;
		fifo[80] <= 0;
		fifo[81] <= 0;
		fifo[82] <= 0;
		fifo[83] <= 0;
		fifo[84] <= 0;
		fifo[85] <= 0;
		fifo[86] <= 0;
		fifo[87] <= 0;
		fifo[88] <= 0;
		fifo[89] <= 0;
		fifo[90] <= 0;
		fifo[91] <= 0;
		fifo[92] <= 0;
		fifo[93] <= 0;
		fifo[94] <= 0;
		fifo[95] <= 0;
		fifo[96] <= 0;
		fifo[97] <= 0;
		fifo[98] <= 0;
		fifo[99] <= 0;
		fifo[100] <= 0;
	end
	else
	begin
			fifo[0] <= in ;
			fifo[1] <= fifo[0];
			fifo[2] <= fifo[1];
			fifo[3] <= fifo[2];
			fifo[4] <= fifo[3];
			fifo[5] <= fifo[4];
			fifo[6] <= fifo[5];
			fifo[7] <= fifo[6];
			fifo[8] <= fifo[7];
			fifo[9] <= fifo[8];
			fifo[10] <= fifo[9];
			fifo[11] <= fifo[10];
			fifo[12] <= fifo[11];
			fifo[13] <= fifo[12];
			fifo[14] <= fifo[13];
			fifo[15] <= fifo[14];
			fifo[16] <= fifo[15];
			fifo[17] <= fifo[16];
			fifo[18] <= fifo[17];
			fifo[19] <= fifo[18];
			fifo[20] <= fifo[19];
			fifo[21] <= fifo[20];
			fifo[22] <= fifo[21];
			fifo[23] <= fifo[22];
			fifo[24] <= fifo[23];
			fifo[25] <= fifo[24];
			fifo[26] <= fifo[25];
			fifo[27] <= fifo[26];
			fifo[28] <= fifo[27];
			fifo[29] <= fifo[28];
			fifo[30] <= fifo[29];
			fifo[31] <= fifo[30];
			fifo[32] <= fifo[31];
			fifo[33] <= fifo[32];
			fifo[34] <= fifo[33];
			fifo[35] <= fifo[34];
			fifo[36] <= fifo[35];
			fifo[37] <= fifo[36];
			fifo[38] <= fifo[37];
			fifo[39] <= fifo[38];
			fifo[40] <= fifo[39];
			fifo[41] <= fifo[40];
			fifo[42] <= fifo[41];
			fifo[43] <= fifo[42];
			fifo[44] <= fifo[43];
			fifo[45] <= fifo[44];
			fifo[46] <= fifo[45];
			fifo[47] <= fifo[46];
			fifo[48] <= fifo[47];
			fifo[49] <= fifo[48];
			fifo[50] <= fifo[49];
			fifo[51] <= fifo[50];
			fifo[52] <= fifo[51];
			fifo[53] <= fifo[52];
			fifo[54] <= fifo[53];
			fifo[55] <= fifo[54];
			fifo[56] <= fifo[55];
			fifo[57] <= fifo[56];
			fifo[58] <= fifo[57];
			fifo[59] <= fifo[58];
			fifo[60] <= fifo[59];
			fifo[61] <= fifo[60];
			fifo[62] <= fifo[61];
			fifo[63] <= fifo[62];
			fifo[64] <= fifo[63];
			fifo[65] <= fifo[64];
			fifo[66] <= fifo[65];
			fifo[67] <= fifo[66];
			fifo[68] <= fifo[67];
			fifo[69] <= fifo[68];
			fifo[70] <= fifo[69];
			fifo[71] <= fifo[70];
			fifo[72] <= fifo[71];
			fifo[73] <= fifo[72];
			fifo[74] <= fifo[73];
			fifo[75] <= fifo[74];
			fifo[76] <= fifo[75];
			fifo[77] <= fifo[76];
			fifo[78] <= fifo[77];
			fifo[79] <= fifo[78];
			fifo[80] <= fifo[79];
			fifo[81] <= fifo[80];
			fifo[82] <= fifo[81];
			fifo[83] <= fifo[82];
			fifo[84] <= fifo[83];
			fifo[85] <= fifo[84];
			fifo[86] <= fifo[85];
			fifo[87] <= fifo[86];
			fifo[88] <= fifo[87];
			fifo[89] <= fifo[88];
			fifo[90] <= fifo[89];
			fifo[91] <= fifo[90];
			fifo[92] <= fifo[91];
			fifo[93] <= fifo[92];
			fifo[94] <= fifo[93];
			fifo[95] <= fifo[94];
			fifo[96] <= fifo[95];
			fifo[97] <= fifo[96];
			fifo[98] <= fifo[97];
			fifo[99] <= fifo[98];
			fifo[100] <= fifo[99];
	end
end

endmodule