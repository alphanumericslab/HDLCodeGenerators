`timescale 1ns / 1ps

module MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL
#(
parameter IN_WIDTH = 16,
parameter INPUT_REG_DEPTH = 1,
parameter MULT_PIPE_DEPTH = 1
)(
input clk, reset, enable,
output reg rowSetInNo = 0,
input inReady,
input signed [IN_WIDTH-1:0] AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
input signed [IN_WIDTH-1:0] AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
input signed [IN_WIDTH-1:0] AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
input signed [IN_WIDTH-1:0] AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
input signed [IN_WIDTH-1:0] AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
input signed [IN_WIDTH-1:0] AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
input signed [IN_WIDTH-1:0] AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
input signed [IN_WIDTH-1:0] AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
input signed [IN_WIDTH-1:0] AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
input signed [IN_WIDTH-1:0] AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
input signed [IN_WIDTH-1:0] VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
output E0toE9Ready,
output reg NUCReady = 0, //not used
output reg rowSetOutNo = 0,
output signed [(2*IN_WIDTH)+3:0] E0, E1, E2, E3, E4, E5, E6, E7, E8, E9, 
output earlyE0toE9Ready,
output reg NUearlyCReady = 0 //not used
);


DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_0 (clk, reset, enable,
inReady,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
E0toE9Ready,
E0,
earlyE0toE9Ready
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_1 (clk, reset, enable,
inReady,
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady1, //not used
E1,
DPearlyOutReady1 //not used
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_2 (clk, reset, enable,
inReady,
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady2, //not used
E2,
DPearlyOutReady2 //not used
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_3 (clk, reset, enable,
inReady,
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady3, //not used
E3,
DPearlyOutReady3 //not used
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_4 (clk, reset, enable,
inReady,
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady4, //not used
E4,
DPearlyOutReady4 //not used
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_5 (clk, reset, enable,
inReady,
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady5, //not used
E5,
DPearlyOutReady5 //not used
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_6 (clk, reset, enable,
inReady,
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady6, //not used
E6,
DPearlyOutReady6 //not used
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_7 (clk, reset, enable,
inReady,
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady7, //not used
E7,
DPearlyOutReady7 //not used
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_8 (clk, reset, enable,
inReady,
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady8, //not used
E8,
DPearlyOutReady8 //not used
);

DotProduct_Systolic_12
#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
DP_9 (clk, reset, enable,
inReady,
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
VE0, VE1, VE2, VE3, VE4, VE5, VE6, VE7, VE8, VE9, VE10, VE11, 
DPOutReady9, //not used
E9,
DPearlyOutReady9 //not used
);

endmodule
