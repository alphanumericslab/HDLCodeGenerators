`ifndef _my_include_vh_
`define _my_include_vh_

`define W 101
`define LOG_W 7
`define DATA_LENGTH  16
`endif
