`timescale 1ns / 1ps

module MatrixAdd_12_10_12PV_noHR_NIR_AXIStream
#(
parameter IN_DATA_LENGHT= 3840, 
parameter OUT_DATA_LENGHT= 2040 
)( 

input aclk,
input aresetn,
input enable,
input [IN_DATA_LENGHT-1:0]s_axi_data,
input s_axi_valid,
input m_axi_ready,
output reg[OUT_DATA_LENGHT-1:0]m_axi_data,
output reg m_axi_valid,
output reg s_axi_ready
);

reg inready;
reg [IN_DATA_LENGHT-1:0]indata;
wire outready;
wire earlyoutready;
wire [OUT_DATA_LENGHT-1:0]outdata;
////////////////instancing wrapping module///////////////////
MatrixAdd_12_10_12PV_noHR_NIR MatrixAdd_12_10_12PV_noHR_NIR_inst(
.clk(aclk),
.reset(!aresetn),
.enable(enable),
.inReady(inready),
.A0V0(indata[3839:3824]),
.A0V1(indata[3839:3824]),
.A0V2(indata[3839:3824]),
.A0V3(indata[3839:3824]),
.A0V4(indata[3839:3824]),
.A0V5(indata[3839:3824]),
.A0V6(indata[3839:3824]),
.A0V7(indata[3839:3824]),
.A0V8(indata[3839:3824]),
.A0V9(indata[3839:3824]),
.A0V10(indata[3839:3824]),
.A0V11(indata[3839:3824]),
.A1V0(indata[3823:3808]),
.A1V1(indata[3823:3808]),
.A1V2(indata[3823:3808]),
.A1V3(indata[3823:3808]),
.A1V4(indata[3823:3808]),
.A1V5(indata[3823:3808]),
.A1V6(indata[3823:3808]),
.A1V7(indata[3823:3808]),
.A1V8(indata[3823:3808]),
.A1V9(indata[3823:3808]),
.A1V10(indata[3823:3808]),
.A1V11(indata[3823:3808]),
.A2V0(indata[3807:3792]),
.A2V1(indata[3807:3792]),
.A2V2(indata[3807:3792]),
.A2V3(indata[3807:3792]),
.A2V4(indata[3807:3792]),
.A2V5(indata[3807:3792]),
.A2V6(indata[3807:3792]),
.A2V7(indata[3807:3792]),
.A2V8(indata[3807:3792]),
.A2V9(indata[3807:3792]),
.A2V10(indata[3807:3792]),
.A2V11(indata[3807:3792]),
.A3V0(indata[3791:3776]),
.A3V1(indata[3791:3776]),
.A3V2(indata[3791:3776]),
.A3V3(indata[3791:3776]),
.A3V4(indata[3791:3776]),
.A3V5(indata[3791:3776]),
.A3V6(indata[3791:3776]),
.A3V7(indata[3791:3776]),
.A3V8(indata[3791:3776]),
.A3V9(indata[3791:3776]),
.A3V10(indata[3791:3776]),
.A3V11(indata[3791:3776]),
.A4V0(indata[3775:3760]),
.A4V1(indata[3775:3760]),
.A4V2(indata[3775:3760]),
.A4V3(indata[3775:3760]),
.A4V4(indata[3775:3760]),
.A4V5(indata[3775:3760]),
.A4V6(indata[3775:3760]),
.A4V7(indata[3775:3760]),
.A4V8(indata[3775:3760]),
.A4V9(indata[3775:3760]),
.A4V10(indata[3775:3760]),
.A4V11(indata[3775:3760]),
.A5V0(indata[3759:3744]),
.A5V1(indata[3759:3744]),
.A5V2(indata[3759:3744]),
.A5V3(indata[3759:3744]),
.A5V4(indata[3759:3744]),
.A5V5(indata[3759:3744]),
.A5V6(indata[3759:3744]),
.A5V7(indata[3759:3744]),
.A5V8(indata[3759:3744]),
.A5V9(indata[3759:3744]),
.A5V10(indata[3759:3744]),
.A5V11(indata[3759:3744]),
.A6V0(indata[3743:3728]),
.A6V1(indata[3743:3728]),
.A6V2(indata[3743:3728]),
.A6V3(indata[3743:3728]),
.A6V4(indata[3743:3728]),
.A6V5(indata[3743:3728]),
.A6V6(indata[3743:3728]),
.A6V7(indata[3743:3728]),
.A6V8(indata[3743:3728]),
.A6V9(indata[3743:3728]),
.A6V10(indata[3743:3728]),
.A6V11(indata[3743:3728]),
.A7V0(indata[3727:3712]),
.A7V1(indata[3727:3712]),
.A7V2(indata[3727:3712]),
.A7V3(indata[3727:3712]),
.A7V4(indata[3727:3712]),
.A7V5(indata[3727:3712]),
.A7V6(indata[3727:3712]),
.A7V7(indata[3727:3712]),
.A7V8(indata[3727:3712]),
.A7V9(indata[3727:3712]),
.A7V10(indata[3727:3712]),
.A7V11(indata[3727:3712]),
.A8V0(indata[3711:3696]),
.A8V1(indata[3711:3696]),
.A8V2(indata[3711:3696]),
.A8V3(indata[3711:3696]),
.A8V4(indata[3711:3696]),
.A8V5(indata[3711:3696]),
.A8V6(indata[3711:3696]),
.A8V7(indata[3711:3696]),
.A8V8(indata[3711:3696]),
.A8V9(indata[3711:3696]),
.A8V10(indata[3711:3696]),
.A8V11(indata[3711:3696]),
.A9V0(indata[3695:3680]),
.A9V1(indata[3695:3680]),
.A9V2(indata[3695:3680]),
.A9V3(indata[3695:3680]),
.A9V4(indata[3695:3680]),
.A9V5(indata[3695:3680]),
.A9V6(indata[3695:3680]),
.A9V7(indata[3695:3680]),
.A9V8(indata[3695:3680]),
.A9V9(indata[3695:3680]),
.A9V10(indata[3695:3680]),
.A9V11(indata[3695:3680]),
.B0V0(indata[1919:1904]),
.B0V1(indata[1919:1904]),
.B0V2(indata[1919:1904]),
.B0V3(indata[1919:1904]),
.B0V4(indata[1919:1904]),
.B0V5(indata[1919:1904]),
.B0V6(indata[1919:1904]),
.B0V7(indata[1919:1904]),
.B0V8(indata[1919:1904]),
.B0V9(indata[1919:1904]),
.B0V10(indata[1919:1904]),
.B0V11(indata[1919:1904]),
.B1V0(indata[1903:1888]),
.B1V1(indata[1903:1888]),
.B1V2(indata[1903:1888]),
.B1V3(indata[1903:1888]),
.B1V4(indata[1903:1888]),
.B1V5(indata[1903:1888]),
.B1V6(indata[1903:1888]),
.B1V7(indata[1903:1888]),
.B1V8(indata[1903:1888]),
.B1V9(indata[1903:1888]),
.B1V10(indata[1903:1888]),
.B1V11(indata[1903:1888]),
.B2V0(indata[1887:1872]),
.B2V1(indata[1887:1872]),
.B2V2(indata[1887:1872]),
.B2V3(indata[1887:1872]),
.B2V4(indata[1887:1872]),
.B2V5(indata[1887:1872]),
.B2V6(indata[1887:1872]),
.B2V7(indata[1887:1872]),
.B2V8(indata[1887:1872]),
.B2V9(indata[1887:1872]),
.B2V10(indata[1887:1872]),
.B2V11(indata[1887:1872]),
.B3V0(indata[1871:1856]),
.B3V1(indata[1871:1856]),
.B3V2(indata[1871:1856]),
.B3V3(indata[1871:1856]),
.B3V4(indata[1871:1856]),
.B3V5(indata[1871:1856]),
.B3V6(indata[1871:1856]),
.B3V7(indata[1871:1856]),
.B3V8(indata[1871:1856]),
.B3V9(indata[1871:1856]),
.B3V10(indata[1871:1856]),
.B3V11(indata[1871:1856]),
.B4V0(indata[1855:1840]),
.B4V1(indata[1855:1840]),
.B4V2(indata[1855:1840]),
.B4V3(indata[1855:1840]),
.B4V4(indata[1855:1840]),
.B4V5(indata[1855:1840]),
.B4V6(indata[1855:1840]),
.B4V7(indata[1855:1840]),
.B4V8(indata[1855:1840]),
.B4V9(indata[1855:1840]),
.B4V10(indata[1855:1840]),
.B4V11(indata[1855:1840]),
.B5V0(indata[1839:1824]),
.B5V1(indata[1839:1824]),
.B5V2(indata[1839:1824]),
.B5V3(indata[1839:1824]),
.B5V4(indata[1839:1824]),
.B5V5(indata[1839:1824]),
.B5V6(indata[1839:1824]),
.B5V7(indata[1839:1824]),
.B5V8(indata[1839:1824]),
.B5V9(indata[1839:1824]),
.B5V10(indata[1839:1824]),
.B5V11(indata[1839:1824]),
.B6V0(indata[1823:1808]),
.B6V1(indata[1823:1808]),
.B6V2(indata[1823:1808]),
.B6V3(indata[1823:1808]),
.B6V4(indata[1823:1808]),
.B6V5(indata[1823:1808]),
.B6V6(indata[1823:1808]),
.B6V7(indata[1823:1808]),
.B6V8(indata[1823:1808]),
.B6V9(indata[1823:1808]),
.B6V10(indata[1823:1808]),
.B6V11(indata[1823:1808]),
.B7V0(indata[1807:1792]),
.B7V1(indata[1807:1792]),
.B7V2(indata[1807:1792]),
.B7V3(indata[1807:1792]),
.B7V4(indata[1807:1792]),
.B7V5(indata[1807:1792]),
.B7V6(indata[1807:1792]),
.B7V7(indata[1807:1792]),
.B7V8(indata[1807:1792]),
.B7V9(indata[1807:1792]),
.B7V10(indata[1807:1792]),
.B7V11(indata[1807:1792]),
.B8V0(indata[1791:1776]),
.B8V1(indata[1791:1776]),
.B8V2(indata[1791:1776]),
.B8V3(indata[1791:1776]),
.B8V4(indata[1791:1776]),
.B8V5(indata[1791:1776]),
.B8V6(indata[1791:1776]),
.B8V7(indata[1791:1776]),
.B8V8(indata[1791:1776]),
.B8V9(indata[1791:1776]),
.B8V10(indata[1791:1776]),
.B8V11(indata[1791:1776]),
.B9V0(indata[1775:1760]),
.B9V1(indata[1775:1760]),
.B9V2(indata[1775:1760]),
.B9V3(indata[1775:1760]),
.B9V4(indata[1775:1760]),
.B9V5(indata[1775:1760]),
.B9V6(indata[1775:1760]),
.B9V7(indata[1775:1760]),
.B9V8(indata[1775:1760]),
.B9V9(indata[1775:1760]),
.B9V10(indata[1775:1760]),
.B9V11(indata[1775:1760]),
.V0toV9outReady(outready),
.S0V0(outdata[2039:2023]),
.S0V1(outdata[2039:2023]),
.S0V2(outdata[2039:2023]),
.S0V3(outdata[2039:2023]),
.S0V4(outdata[2039:2023]),
.S0V5(outdata[2039:2023]),
.S0V6(outdata[2039:2023]),
.S0V7(outdata[2039:2023]),
.S0V8(outdata[2039:2023]),
.S0V9(outdata[2039:2023]),
.S0V10(outdata[2039:2023]),
.S0V11(outdata[2039:2023]),
.S1V0(outdata[2022:2006]),
.S1V1(outdata[2022:2006]),
.S1V2(outdata[2022:2006]),
.S1V3(outdata[2022:2006]),
.S1V4(outdata[2022:2006]),
.S1V5(outdata[2022:2006]),
.S1V6(outdata[2022:2006]),
.S1V7(outdata[2022:2006]),
.S1V8(outdata[2022:2006]),
.S1V9(outdata[2022:2006]),
.S1V10(outdata[2022:2006]),
.S1V11(outdata[2022:2006]),
.S2V0(outdata[2005:1989]),
.S2V1(outdata[2005:1989]),
.S2V2(outdata[2005:1989]),
.S2V3(outdata[2005:1989]),
.S2V4(outdata[2005:1989]),
.S2V5(outdata[2005:1989]),
.S2V6(outdata[2005:1989]),
.S2V7(outdata[2005:1989]),
.S2V8(outdata[2005:1989]),
.S2V9(outdata[2005:1989]),
.S2V10(outdata[2005:1989]),
.S2V11(outdata[2005:1989]),
.S3V0(outdata[1988:1972]),
.S3V1(outdata[1988:1972]),
.S3V2(outdata[1988:1972]),
.S3V3(outdata[1988:1972]),
.S3V4(outdata[1988:1972]),
.S3V5(outdata[1988:1972]),
.S3V6(outdata[1988:1972]),
.S3V7(outdata[1988:1972]),
.S3V8(outdata[1988:1972]),
.S3V9(outdata[1988:1972]),
.S3V10(outdata[1988:1972]),
.S3V11(outdata[1988:1972]),
.S4V0(outdata[1971:1955]),
.S4V1(outdata[1971:1955]),
.S4V2(outdata[1971:1955]),
.S4V3(outdata[1971:1955]),
.S4V4(outdata[1971:1955]),
.S4V5(outdata[1971:1955]),
.S4V6(outdata[1971:1955]),
.S4V7(outdata[1971:1955]),
.S4V8(outdata[1971:1955]),
.S4V9(outdata[1971:1955]),
.S4V10(outdata[1971:1955]),
.S4V11(outdata[1971:1955]),
.S5V0(outdata[1954:1938]),
.S5V1(outdata[1954:1938]),
.S5V2(outdata[1954:1938]),
.S5V3(outdata[1954:1938]),
.S5V4(outdata[1954:1938]),
.S5V5(outdata[1954:1938]),
.S5V6(outdata[1954:1938]),
.S5V7(outdata[1954:1938]),
.S5V8(outdata[1954:1938]),
.S5V9(outdata[1954:1938]),
.S5V10(outdata[1954:1938]),
.S5V11(outdata[1954:1938]),
.S6V0(outdata[1937:1921]),
.S6V1(outdata[1937:1921]),
.S6V2(outdata[1937:1921]),
.S6V3(outdata[1937:1921]),
.S6V4(outdata[1937:1921]),
.S6V5(outdata[1937:1921]),
.S6V6(outdata[1937:1921]),
.S6V7(outdata[1937:1921]),
.S6V8(outdata[1937:1921]),
.S6V9(outdata[1937:1921]),
.S6V10(outdata[1937:1921]),
.S6V11(outdata[1937:1921]),
.S7V0(outdata[1920:1904]),
.S7V1(outdata[1920:1904]),
.S7V2(outdata[1920:1904]),
.S7V3(outdata[1920:1904]),
.S7V4(outdata[1920:1904]),
.S7V5(outdata[1920:1904]),
.S7V6(outdata[1920:1904]),
.S7V7(outdata[1920:1904]),
.S7V8(outdata[1920:1904]),
.S7V9(outdata[1920:1904]),
.S7V10(outdata[1920:1904]),
.S7V11(outdata[1920:1904]),
.S8V0(outdata[1903:1887]),
.S8V1(outdata[1903:1887]),
.S8V2(outdata[1903:1887]),
.S8V3(outdata[1903:1887]),
.S8V4(outdata[1903:1887]),
.S8V5(outdata[1903:1887]),
.S8V6(outdata[1903:1887]),
.S8V7(outdata[1903:1887]),
.S8V8(outdata[1903:1887]),
.S8V9(outdata[1903:1887]),
.S8V10(outdata[1903:1887]),
.S8V11(outdata[1903:1887]),
.S9V0(outdata[1886:1870]),
.S9V1(outdata[1886:1870]),
.S9V2(outdata[1886:1870]),
.S9V3(outdata[1886:1870]),
.S9V4(outdata[1886:1870]),
.S9V5(outdata[1886:1870]),
.S9V6(outdata[1886:1870]),
.S9V7(outdata[1886:1870]),
.S9V8(outdata[1886:1870]),
.S9V9(outdata[1886:1870]),
.S9V10(outdata[1886:1870]),
.S9V11(outdata[1886:1870]),
.V0toV10earlyOutReady(earlyoutready)
);
/////////////////Main body/////////////
always @(posedge aclk)begin
 if(aresetn==0)begin
  m_axi_data<=0;
  m_axi_valid<=0;
 end
 else begin
  if(m_axi_ready==1 && m_axi_valid==1)begin
   m_axi_valid<=0;
  end
  else if(outready==1)begin
   m_axi_valid<=1;
   m_axi_data<=outdata;
  end
 end
end
always @(posedge aclk)begin
 if(aresetn==0)begin
  s_axi_ready<=1;
  inready<=0;
  indata<=0;
 end
 else begin
  inready<=0;
  if(s_axi_valid==1 && s_axi_ready==1)begin
   s_axi_ready<=0;
   inready<=1;
   indata<= s_axi_data;
  end
  else if(m_axi_valid==1 && m_axi_ready==1)begin
   s_axi_ready<=1;
  end
 end
end

endmodule
