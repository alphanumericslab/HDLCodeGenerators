`timescale 1ns / 1ps

module MatrixMatrixMultiply_10_12_10_10PR_10PC_noHR_C12_A0_NCL_NRL.v
#(
parameter IN_WIDTH = 16,
parameter INPUT_REG_DEPTH = 1,
parameter MULT_PIPE_DEPTH = 1
)(
input clk, reset, enable,
output rowSetInNo,
output reg columnSetInNo = 0,
input inReady,
input signed [IN_WIDTH-1:0] AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
input signed [IN_WIDTH-1:0] BE0C0, BE1C0, BE2C0, BE3C0, BE4C0, BE5C0, BE6C0, BE7C0, BE8C0, BE9C0, BE10C0, BE11C0, 
BE0C1, BE1C1, BE2C1, BE3C1, BE4C1, BE5C1, BE6C1, BE7C1, BE8C1, BE9C1, BE10C1, BE11C1, 
BE0C2, BE1C2, BE2C2, BE3C2, BE4C2, BE5C2, BE6C2, BE7C2, BE8C2, BE9C2, BE10C2, BE11C2, 
BE0C3, BE1C3, BE2C3, BE3C3, BE4C3, BE5C3, BE6C3, BE7C3, BE8C3, BE9C3, BE10C3, BE11C3, 
BE0C4, BE1C4, BE2C4, BE3C4, BE4C4, BE5C4, BE6C4, BE7C4, BE8C4, BE9C4, BE10C4, BE11C4, 
BE0C5, BE1C5, BE2C5, BE3C5, BE4C5, BE5C5, BE6C5, BE7C5, BE8C5, BE9C5, BE10C5, BE11C5, 
BE0C6, BE1C6, BE2C6, BE3C6, BE4C6, BE5C6, BE6C6, BE7C6, BE8C6, BE9C6, BE10C6, BE11C6, 
BE0C7, BE1C7, BE2C7, BE3C7, BE4C7, BE5C7, BE6C7, BE7C7, BE8C7, BE9C7, BE10C7, BE11C7, 
BE0C8, BE1C8, BE2C8, BE3C8, BE4C8, BE5C8, BE6C8, BE7C8, BE8C8, BE9C8, BE10C8, BE11C8, 
BE0C9, BE1C9, BE2C9, BE3C9, BE4C9, BE5C9, BE6C9, BE7C9, BE8C9, BE9C9, BE10C9, BE11C9, 
output C0toC9R0toR9EReady,
output reg NUEReady1 = 0, //not used
output reg NUEReady2 = 0, //not used
output reg NUEReady3 = 0, //not used
output rowSetOutNo,
output reg columnSetOutNo = 0,
output signed [(2*IN_WIDTH)+3:0] EC0R0, EC0R1, EC0R2, EC0R3, EC0R4, EC0R5, EC0R6, EC0R7, EC0R8, EC0R9, EC1R0, EC1R1, EC1R2, EC1R3, EC1R4, EC1R5, EC1R6, EC1R7, EC1R8, EC1R9, EC2R0, EC2R1, EC2R2, EC2R3, EC2R4, EC2R5, EC2R6, EC2R7, EC2R8, EC2R9, EC3R0, EC3R1, EC3R2, EC3R3, EC3R4, EC3R5, EC3R6, EC3R7, EC3R8, EC3R9, EC4R0, EC4R1, EC4R2, EC4R3, EC4R4, EC4R5, EC4R6, EC4R7, EC4R8, EC4R9, EC5R0, EC5R1, EC5R2, EC5R3, EC5R4, EC5R5, EC5R6, EC5R7, EC5R8, EC5R9, EC6R0, EC6R1, EC6R2, EC6R3, EC6R4, EC6R5, EC6R6, EC6R7, EC6R8, EC6R9, EC7R0, EC7R1, EC7R2, EC7R3, EC7R4, EC7R5, EC7R6, EC7R7, EC7R8, EC7R9, EC8R0, EC8R1, EC8R2, EC8R3, EC8R4, EC8R5, EC8R6, EC8R7, EC8R8, EC8R9, EC9R0, EC9R1, EC9R2, EC9R3, EC9R4, EC9R5, EC9R6, EC9R7, EC9R8, EC9R9, 
output earlyC0toC9R0toR9EReady,
output reg NUeEReady1 = 0, //not used
output reg NUeEReady2 = 0, //not used
output reg NUeEReady3 = 0 //not used
);

wire inReadyC = inReady;
wire gettingIn = 1; //for simulation
MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_0(clk, reset, enable,
rowSetInNo,
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C0, BE1C0, BE2C0, BE3C0, BE4C0, BE5C0, BE6C0, BE7C0, BE8C0, BE9C0, BE10C0, BE11C0, 
C0toC9R0toR9EReady,
LLMVMoutReadyA0, //not used
rowSetOutNo,
EC0R0,
EC0R1,
EC0R2,
EC0R3,
EC0R4,
EC0R5,
EC0R6,
EC0R7,
EC0R8,
EC0R9,
earlyC0toC9R0toR9EReady,
LLMVMearlyOutReadyA0 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_1(clk, reset, enable,
LLrowSetInNo1, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C1, BE1C1, BE2C1, BE3C1, BE4C1, BE5C1, BE6C1, BE7C1, BE8C1, BE9C1, BE10C1, BE11C1, 
LLMVMoutReady1, //not used
LLMVMoutReadyA1, //not used
LLrowSetOutNo1, //not used
EC1R0,
EC1R1,
EC1R2,
EC1R3,
EC1R4,
EC1R5,
EC1R6,
EC1R7,
EC1R8,
EC1R9,
LLMVMearlyOutReady1,
LLMVMearlyOutReadyA1 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_2(clk, reset, enable,
LLrowSetInNo2, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C2, BE1C2, BE2C2, BE3C2, BE4C2, BE5C2, BE6C2, BE7C2, BE8C2, BE9C2, BE10C2, BE11C2, 
LLMVMoutReady2, //not used
LLMVMoutReadyA2, //not used
LLrowSetOutNo2, //not used
EC2R0,
EC2R1,
EC2R2,
EC2R3,
EC2R4,
EC2R5,
EC2R6,
EC2R7,
EC2R8,
EC2R9,
LLMVMearlyOutReady2,
LLMVMearlyOutReadyA2 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_3(clk, reset, enable,
LLrowSetInNo3, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C3, BE1C3, BE2C3, BE3C3, BE4C3, BE5C3, BE6C3, BE7C3, BE8C3, BE9C3, BE10C3, BE11C3, 
LLMVMoutReady3, //not used
LLMVMoutReadyA3, //not used
LLrowSetOutNo3, //not used
EC3R0,
EC3R1,
EC3R2,
EC3R3,
EC3R4,
EC3R5,
EC3R6,
EC3R7,
EC3R8,
EC3R9,
LLMVMearlyOutReady3,
LLMVMearlyOutReadyA3 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_4(clk, reset, enable,
LLrowSetInNo4, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C4, BE1C4, BE2C4, BE3C4, BE4C4, BE5C4, BE6C4, BE7C4, BE8C4, BE9C4, BE10C4, BE11C4, 
LLMVMoutReady4, //not used
LLMVMoutReadyA4, //not used
LLrowSetOutNo4, //not used
EC4R0,
EC4R1,
EC4R2,
EC4R3,
EC4R4,
EC4R5,
EC4R6,
EC4R7,
EC4R8,
EC4R9,
LLMVMearlyOutReady4,
LLMVMearlyOutReadyA4 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_5(clk, reset, enable,
LLrowSetInNo5, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C5, BE1C5, BE2C5, BE3C5, BE4C5, BE5C5, BE6C5, BE7C5, BE8C5, BE9C5, BE10C5, BE11C5, 
LLMVMoutReady5, //not used
LLMVMoutReadyA5, //not used
LLrowSetOutNo5, //not used
EC5R0,
EC5R1,
EC5R2,
EC5R3,
EC5R4,
EC5R5,
EC5R6,
EC5R7,
EC5R8,
EC5R9,
LLMVMearlyOutReady5,
LLMVMearlyOutReadyA5 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_6(clk, reset, enable,
LLrowSetInNo6, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C6, BE1C6, BE2C6, BE3C6, BE4C6, BE5C6, BE6C6, BE7C6, BE8C6, BE9C6, BE10C6, BE11C6, 
LLMVMoutReady6, //not used
LLMVMoutReadyA6, //not used
LLrowSetOutNo6, //not used
EC6R0,
EC6R1,
EC6R2,
EC6R3,
EC6R4,
EC6R5,
EC6R6,
EC6R7,
EC6R8,
EC6R9,
LLMVMearlyOutReady6,
LLMVMearlyOutReadyA6 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_7(clk, reset, enable,
LLrowSetInNo7, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C7, BE1C7, BE2C7, BE3C7, BE4C7, BE5C7, BE6C7, BE7C7, BE8C7, BE9C7, BE10C7, BE11C7, 
LLMVMoutReady7, //not used
LLMVMoutReadyA7, //not used
LLrowSetOutNo7, //not used
EC7R0,
EC7R1,
EC7R2,
EC7R3,
EC7R4,
EC7R5,
EC7R6,
EC7R7,
EC7R8,
EC7R9,
LLMVMearlyOutReady7,
LLMVMearlyOutReadyA7 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_8(clk, reset, enable,
LLrowSetInNo8, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C8, BE1C8, BE2C8, BE3C8, BE4C8, BE5C8, BE6C8, BE7C8, BE8C8, BE9C8, BE10C8, BE11C8, 
LLMVMoutReady8, //not used
LLMVMoutReadyA8, //not used
LLrowSetOutNo8, //not used
EC8R0,
EC8R1,
EC8R2,
EC8R3,
EC8R4,
EC8R5,
EC8R6,
EC8R7,
EC8R8,
EC8R9,
LLMVMearlyOutReady8,
LLMVMearlyOutReadyA8 //not used
);

MatrixVectorMultiply_10_12_10PR_noHR_C12_A0_NVL#( .IN_WIDTH(IN_WIDTH), .INPUT_REG_DEPTH(INPUT_REG_DEPTH), .MULT_PIPE_DEPTH(MULT_PIPE_DEPTH) )
MVM_9(clk, reset, enable,
LLrowSetInNo9, //not used
inReadyC,
AE0R0, AE1R0, AE2R0, AE3R0, AE4R0, AE5R0, AE6R0, AE7R0, AE8R0, AE9R0, AE10R0, AE11R0, 
AE0R1, AE1R1, AE2R1, AE3R1, AE4R1, AE5R1, AE6R1, AE7R1, AE8R1, AE9R1, AE10R1, AE11R1, 
AE0R2, AE1R2, AE2R2, AE3R2, AE4R2, AE5R2, AE6R2, AE7R2, AE8R2, AE9R2, AE10R2, AE11R2, 
AE0R3, AE1R3, AE2R3, AE3R3, AE4R3, AE5R3, AE6R3, AE7R3, AE8R3, AE9R3, AE10R3, AE11R3, 
AE0R4, AE1R4, AE2R4, AE3R4, AE4R4, AE5R4, AE6R4, AE7R4, AE8R4, AE9R4, AE10R4, AE11R4, 
AE0R5, AE1R5, AE2R5, AE3R5, AE4R5, AE5R5, AE6R5, AE7R5, AE8R5, AE9R5, AE10R5, AE11R5, 
AE0R6, AE1R6, AE2R6, AE3R6, AE4R6, AE5R6, AE6R6, AE7R6, AE8R6, AE9R6, AE10R6, AE11R6, 
AE0R7, AE1R7, AE2R7, AE3R7, AE4R7, AE5R7, AE6R7, AE7R7, AE8R7, AE9R7, AE10R7, AE11R7, 
AE0R8, AE1R8, AE2R8, AE3R8, AE4R8, AE5R8, AE6R8, AE7R8, AE8R8, AE9R8, AE10R8, AE11R8, 
AE0R9, AE1R9, AE2R9, AE3R9, AE4R9, AE5R9, AE6R9, AE7R9, AE8R9, AE9R9, AE10R9, AE11R9, 
BE0C9, BE1C9, BE2C9, BE3C9, BE4C9, BE5C9, BE6C9, BE7C9, BE8C9, BE9C9, BE10C9, BE11C9, 
LLMVMoutReady9, //not used
LLMVMoutReadyA9, //not used
LLrowSetOutNo9, //not used
EC9R0,
EC9R1,
EC9R2,
EC9R3,
EC9R4,
EC9R5,
EC9R6,
EC9R7,
EC9R8,
EC9R9,
LLMVMearlyOutReady9,
LLMVMearlyOutReadyA9 //not used
);

endmodule
