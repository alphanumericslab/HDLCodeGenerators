`timescale 1ns / 1ps
`include "macro.vh"
///////////////////////
module top ( clk ,reset ,X ,median );

output [`DATA_LENGTH-1:0] median ;
input [`DATA_LENGTH-1:0] X ;
input clk ,reset ;

wire 	[`DATA_LENGTH-1:0] R_old, R1 ,R2 ,R3 ,R4 ,R5 ,R6 ,R7 ,R8 ,R9 ,R10 ,R11 ,R12 ,R13 ,R14 ,R15 ,R16 ,R17 ,R18 ,R19 ,R20 ,R21 ,R22 ,R23 ,R24 ,R25 ,R26 ,R27 ,R28 ,R29 ,R30 ,R31 ,R32 ,R33 ,R34 ,R35 ,R36 ,R37 ,R38 ,R39 ,R40 ,R41 ,R42 ,R43 ,R44 ,R45 ,R46 ,R47 ,R48 ,R49 ,R50 ,R51 ,R52 ,R53 ,R54 ,R55 ,R56 ,R57 ,R58 ,R59 ,R60 ,R61 ,R62 ,R63 ,R64 ,R65 ,R66 ,R67 ,R68 ,R69 ,R70 ,R71 ,R72 ,R73 ,R74 ,R75 ,R76 ,R77 ,R78 ,R79 ,R80 ,R81 ,R82 ,R83 ,R84 ,R85 ,R86 ,R87 ,R88 ,R89 ,R90 ,R91 ,R92 ,R93 ,R94 ,R95 ,R96 ,R97 ,R98 ,R99 ,R100 ,R101;
wire 	T1 ,T2 ,T3 ,T4 ,T5 ,T6 ,T7 ,T8 ,T9 ,T10 ,T11 ,T12 ,T13 ,T14 ,T15 ,T16 ,T17 ,T18 ,T19 ,T20 ,T21 ,T22 ,T23 ,T24 ,T25 ,T26 ,T27 ,T28 ,T29 ,T30 ,T31 ,T32 ,T33 ,T34 ,T35 ,T36 ,T37 ,T38 ,T39 ,T40 ,T41 ,T42 ,T43 ,T44 ,T45 ,T46 ,T47 ,T48 ,T49 ,T50 ,T51 ,T52 ,T53 ,T54 ,T55 ,T56 ,T57 ,T58 ,T59 ,T60 ,T61 ,T62 ,T63 ,T64 ,T65 ,T66 ,T67 ,T68 ,T69 ,T70 ,T71 ,T72 ,T73 ,T74 ,T75 ,T76 ,T77 ,T78 ,T79 ,T80 ,T81 ,T82 ,T83 ,T84 ,T85 ,T86 ,T87 ,T88 ,T89 ,T90 ,T91 ,T92 ,T93 ,T94 ,T95 ,T96 ,T97 ,T98 ,T99 ,T100 ,T101;
wire 	 Z1 ,Z2 ,Z3 ,Z4 ,Z5 ,Z6 ,Z7 ,Z8 ,Z9 ,Z10 ,Z11 ,Z12 ,Z13 ,Z14 ,Z15 ,Z16 ,Z17 ,Z18 ,Z19 ,Z20 ,Z21 ,Z22 ,Z23 ,Z24 ,Z25 ,Z26 ,Z27 ,Z28 ,Z29 ,Z30 ,Z31 ,Z32 ,Z33 ,Z34 ,Z35 ,Z36 ,Z37 ,Z38 ,Z39 ,Z40 ,Z41 ,Z42 ,Z43 ,Z44 ,Z45 ,Z46 ,Z47 ,Z48 ,Z49 ,Z50 ,Z51 ,Z52 ,Z53 ,Z54 ,Z55 ,Z56 ,Z57 ,Z58 ,Z59 ,Z60 ,Z61 ,Z62 ,Z63 ,Z64 ,Z65 ,Z66 ,Z67 ,Z68 ,Z69 ,Z70 ,Z71 ,Z72 ,Z73 ,Z74 ,Z75 ,Z76 ,Z77 ,Z78 ,Z79 ,Z80 ,Z81 ,Z82 ,Z83 ,Z84 ,Z85 ,Z86 ,Z87 ,Z88 ,Z89 ,Z90 ,Z91 ,Z92 ,Z93 ,Z94 ,Z95 ,Z96 ,Z97 ,Z98 ,Z99 ,Z100;
assign median =  R51;

FIFO myfifo(.in(X), .out(R_old), .clk(clk), .reset(reset));
medianCell_leftMst  m1(.X(X) , .clk(clk), .reset(reset) , .R_R(R2), .T_R(T2), .R_old(R_old), .Z(Z1), .R(R1), .T(T1));
medianFilterCell  m2(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z1), .R_L(R1),.R_R(R3) ,.T_L(T1), .T_R(T3), .R_old(R_old), .Z(Z2), .R(R2), .T(T2));
medianFilterCell  m3(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z2), .R_L(R2),.R_R(R4) ,.T_L(T2), .T_R(T4), .R_old(R_old), .Z(Z3), .R(R3), .T(T3));
medianFilterCell  m4(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z3), .R_L(R3),.R_R(R5) ,.T_L(T3), .T_R(T5), .R_old(R_old), .Z(Z4), .R(R4), .T(T4));
medianFilterCell  m5(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z4), .R_L(R4),.R_R(R6) ,.T_L(T4), .T_R(T6), .R_old(R_old), .Z(Z5), .R(R5), .T(T5));
medianFilterCell  m6(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z5), .R_L(R5),.R_R(R7) ,.T_L(T5), .T_R(T7), .R_old(R_old), .Z(Z6), .R(R6), .T(T6));
medianFilterCell  m7(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z6), .R_L(R6),.R_R(R8) ,.T_L(T6), .T_R(T8), .R_old(R_old), .Z(Z7), .R(R7), .T(T7));
medianFilterCell  m8(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z7), .R_L(R7),.R_R(R9) ,.T_L(T7), .T_R(T9), .R_old(R_old), .Z(Z8), .R(R8), .T(T8));
medianFilterCell  m9(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z8), .R_L(R8),.R_R(R10) ,.T_L(T8), .T_R(T10), .R_old(R_old), .Z(Z9), .R(R9), .T(T9));
medianFilterCell  m10(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z9), .R_L(R9),.R_R(R11) ,.T_L(T9), .T_R(T11), .R_old(R_old), .Z(Z10), .R(R10), .T(T10));
medianFilterCell  m11(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z10), .R_L(R10),.R_R(R12) ,.T_L(T10), .T_R(T12), .R_old(R_old), .Z(Z11), .R(R11), .T(T11));
medianFilterCell  m12(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z11), .R_L(R11),.R_R(R13) ,.T_L(T11), .T_R(T13), .R_old(R_old), .Z(Z12), .R(R12), .T(T12));
medianFilterCell  m13(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z12), .R_L(R12),.R_R(R14) ,.T_L(T12), .T_R(T14), .R_old(R_old), .Z(Z13), .R(R13), .T(T13));
medianFilterCell  m14(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z13), .R_L(R13),.R_R(R15) ,.T_L(T13), .T_R(T15), .R_old(R_old), .Z(Z14), .R(R14), .T(T14));
medianFilterCell  m15(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z14), .R_L(R14),.R_R(R16) ,.T_L(T14), .T_R(T16), .R_old(R_old), .Z(Z15), .R(R15), .T(T15));
medianFilterCell  m16(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z15), .R_L(R15),.R_R(R17) ,.T_L(T15), .T_R(T17), .R_old(R_old), .Z(Z16), .R(R16), .T(T16));
medianFilterCell  m17(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z16), .R_L(R16),.R_R(R18) ,.T_L(T16), .T_R(T18), .R_old(R_old), .Z(Z17), .R(R17), .T(T17));
medianFilterCell  m18(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z17), .R_L(R17),.R_R(R19) ,.T_L(T17), .T_R(T19), .R_old(R_old), .Z(Z18), .R(R18), .T(T18));
medianFilterCell  m19(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z18), .R_L(R18),.R_R(R20) ,.T_L(T18), .T_R(T20), .R_old(R_old), .Z(Z19), .R(R19), .T(T19));
medianFilterCell  m20(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z19), .R_L(R19),.R_R(R21) ,.T_L(T19), .T_R(T21), .R_old(R_old), .Z(Z20), .R(R20), .T(T20));
medianFilterCell  m21(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z20), .R_L(R20),.R_R(R22) ,.T_L(T20), .T_R(T22), .R_old(R_old), .Z(Z21), .R(R21), .T(T21));
medianFilterCell  m22(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z21), .R_L(R21),.R_R(R23) ,.T_L(T21), .T_R(T23), .R_old(R_old), .Z(Z22), .R(R22), .T(T22));
medianFilterCell  m23(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z22), .R_L(R22),.R_R(R24) ,.T_L(T22), .T_R(T24), .R_old(R_old), .Z(Z23), .R(R23), .T(T23));
medianFilterCell  m24(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z23), .R_L(R23),.R_R(R25) ,.T_L(T23), .T_R(T25), .R_old(R_old), .Z(Z24), .R(R24), .T(T24));
medianFilterCell  m25(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z24), .R_L(R24),.R_R(R26) ,.T_L(T24), .T_R(T26), .R_old(R_old), .Z(Z25), .R(R25), .T(T25));
medianFilterCell  m26(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z25), .R_L(R25),.R_R(R27) ,.T_L(T25), .T_R(T27), .R_old(R_old), .Z(Z26), .R(R26), .T(T26));
medianFilterCell  m27(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z26), .R_L(R26),.R_R(R28) ,.T_L(T26), .T_R(T28), .R_old(R_old), .Z(Z27), .R(R27), .T(T27));
medianFilterCell  m28(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z27), .R_L(R27),.R_R(R29) ,.T_L(T27), .T_R(T29), .R_old(R_old), .Z(Z28), .R(R28), .T(T28));
medianFilterCell  m29(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z28), .R_L(R28),.R_R(R30) ,.T_L(T28), .T_R(T30), .R_old(R_old), .Z(Z29), .R(R29), .T(T29));
medianFilterCell  m30(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z29), .R_L(R29),.R_R(R31) ,.T_L(T29), .T_R(T31), .R_old(R_old), .Z(Z30), .R(R30), .T(T30));
medianFilterCell  m31(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z30), .R_L(R30),.R_R(R32) ,.T_L(T30), .T_R(T32), .R_old(R_old), .Z(Z31), .R(R31), .T(T31));
medianFilterCell  m32(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z31), .R_L(R31),.R_R(R33) ,.T_L(T31), .T_R(T33), .R_old(R_old), .Z(Z32), .R(R32), .T(T32));
medianFilterCell  m33(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z32), .R_L(R32),.R_R(R34) ,.T_L(T32), .T_R(T34), .R_old(R_old), .Z(Z33), .R(R33), .T(T33));
medianFilterCell  m34(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z33), .R_L(R33),.R_R(R35) ,.T_L(T33), .T_R(T35), .R_old(R_old), .Z(Z34), .R(R34), .T(T34));
medianFilterCell  m35(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z34), .R_L(R34),.R_R(R36) ,.T_L(T34), .T_R(T36), .R_old(R_old), .Z(Z35), .R(R35), .T(T35));
medianFilterCell  m36(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z35), .R_L(R35),.R_R(R37) ,.T_L(T35), .T_R(T37), .R_old(R_old), .Z(Z36), .R(R36), .T(T36));
medianFilterCell  m37(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z36), .R_L(R36),.R_R(R38) ,.T_L(T36), .T_R(T38), .R_old(R_old), .Z(Z37), .R(R37), .T(T37));
medianFilterCell  m38(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z37), .R_L(R37),.R_R(R39) ,.T_L(T37), .T_R(T39), .R_old(R_old), .Z(Z38), .R(R38), .T(T38));
medianFilterCell  m39(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z38), .R_L(R38),.R_R(R40) ,.T_L(T38), .T_R(T40), .R_old(R_old), .Z(Z39), .R(R39), .T(T39));
medianFilterCell  m40(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z39), .R_L(R39),.R_R(R41) ,.T_L(T39), .T_R(T41), .R_old(R_old), .Z(Z40), .R(R40), .T(T40));
medianFilterCell  m41(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z40), .R_L(R40),.R_R(R42) ,.T_L(T40), .T_R(T42), .R_old(R_old), .Z(Z41), .R(R41), .T(T41));
medianFilterCell  m42(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z41), .R_L(R41),.R_R(R43) ,.T_L(T41), .T_R(T43), .R_old(R_old), .Z(Z42), .R(R42), .T(T42));
medianFilterCell  m43(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z42), .R_L(R42),.R_R(R44) ,.T_L(T42), .T_R(T44), .R_old(R_old), .Z(Z43), .R(R43), .T(T43));
medianFilterCell  m44(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z43), .R_L(R43),.R_R(R45) ,.T_L(T43), .T_R(T45), .R_old(R_old), .Z(Z44), .R(R44), .T(T44));
medianFilterCell  m45(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z44), .R_L(R44),.R_R(R46) ,.T_L(T44), .T_R(T46), .R_old(R_old), .Z(Z45), .R(R45), .T(T45));
medianFilterCell  m46(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z45), .R_L(R45),.R_R(R47) ,.T_L(T45), .T_R(T47), .R_old(R_old), .Z(Z46), .R(R46), .T(T46));
medianFilterCell  m47(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z46), .R_L(R46),.R_R(R48) ,.T_L(T46), .T_R(T48), .R_old(R_old), .Z(Z47), .R(R47), .T(T47));
medianFilterCell  m48(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z47), .R_L(R47),.R_R(R49) ,.T_L(T47), .T_R(T49), .R_old(R_old), .Z(Z48), .R(R48), .T(T48));
medianFilterCell  m49(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z48), .R_L(R48),.R_R(R50) ,.T_L(T48), .T_R(T50), .R_old(R_old), .Z(Z49), .R(R49), .T(T49));
medianFilterCell  m50(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z49), .R_L(R49),.R_R(R51) ,.T_L(T49), .T_R(T51), .R_old(R_old), .Z(Z50), .R(R50), .T(T50));
medianFilterCell  m51(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z50), .R_L(R50),.R_R(R52) ,.T_L(T50), .T_R(T52), .R_old(R_old), .Z(Z51), .R(R51), .T(T51));
medianFilterCell  m52(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z51), .R_L(R51),.R_R(R53) ,.T_L(T51), .T_R(T53), .R_old(R_old), .Z(Z52), .R(R52), .T(T52));
medianFilterCell  m53(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z52), .R_L(R52),.R_R(R54) ,.T_L(T52), .T_R(T54), .R_old(R_old), .Z(Z53), .R(R53), .T(T53));
medianFilterCell  m54(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z53), .R_L(R53),.R_R(R55) ,.T_L(T53), .T_R(T55), .R_old(R_old), .Z(Z54), .R(R54), .T(T54));
medianFilterCell  m55(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z54), .R_L(R54),.R_R(R56) ,.T_L(T54), .T_R(T56), .R_old(R_old), .Z(Z55), .R(R55), .T(T55));
medianFilterCell  m56(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z55), .R_L(R55),.R_R(R57) ,.T_L(T55), .T_R(T57), .R_old(R_old), .Z(Z56), .R(R56), .T(T56));
medianFilterCell  m57(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z56), .R_L(R56),.R_R(R58) ,.T_L(T56), .T_R(T58), .R_old(R_old), .Z(Z57), .R(R57), .T(T57));
medianFilterCell  m58(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z57), .R_L(R57),.R_R(R59) ,.T_L(T57), .T_R(T59), .R_old(R_old), .Z(Z58), .R(R58), .T(T58));
medianFilterCell  m59(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z58), .R_L(R58),.R_R(R60) ,.T_L(T58), .T_R(T60), .R_old(R_old), .Z(Z59), .R(R59), .T(T59));
medianFilterCell  m60(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z59), .R_L(R59),.R_R(R61) ,.T_L(T59), .T_R(T61), .R_old(R_old), .Z(Z60), .R(R60), .T(T60));
medianFilterCell  m61(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z60), .R_L(R60),.R_R(R62) ,.T_L(T60), .T_R(T62), .R_old(R_old), .Z(Z61), .R(R61), .T(T61));
medianFilterCell  m62(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z61), .R_L(R61),.R_R(R63) ,.T_L(T61), .T_R(T63), .R_old(R_old), .Z(Z62), .R(R62), .T(T62));
medianFilterCell  m63(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z62), .R_L(R62),.R_R(R64) ,.T_L(T62), .T_R(T64), .R_old(R_old), .Z(Z63), .R(R63), .T(T63));
medianFilterCell  m64(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z63), .R_L(R63),.R_R(R65) ,.T_L(T63), .T_R(T65), .R_old(R_old), .Z(Z64), .R(R64), .T(T64));
medianFilterCell  m65(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z64), .R_L(R64),.R_R(R66) ,.T_L(T64), .T_R(T66), .R_old(R_old), .Z(Z65), .R(R65), .T(T65));
medianFilterCell  m66(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z65), .R_L(R65),.R_R(R67) ,.T_L(T65), .T_R(T67), .R_old(R_old), .Z(Z66), .R(R66), .T(T66));
medianFilterCell  m67(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z66), .R_L(R66),.R_R(R68) ,.T_L(T66), .T_R(T68), .R_old(R_old), .Z(Z67), .R(R67), .T(T67));
medianFilterCell  m68(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z67), .R_L(R67),.R_R(R69) ,.T_L(T67), .T_R(T69), .R_old(R_old), .Z(Z68), .R(R68), .T(T68));
medianFilterCell  m69(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z68), .R_L(R68),.R_R(R70) ,.T_L(T68), .T_R(T70), .R_old(R_old), .Z(Z69), .R(R69), .T(T69));
medianFilterCell  m70(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z69), .R_L(R69),.R_R(R71) ,.T_L(T69), .T_R(T71), .R_old(R_old), .Z(Z70), .R(R70), .T(T70));
medianFilterCell  m71(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z70), .R_L(R70),.R_R(R72) ,.T_L(T70), .T_R(T72), .R_old(R_old), .Z(Z71), .R(R71), .T(T71));
medianFilterCell  m72(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z71), .R_L(R71),.R_R(R73) ,.T_L(T71), .T_R(T73), .R_old(R_old), .Z(Z72), .R(R72), .T(T72));
medianFilterCell  m73(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z72), .R_L(R72),.R_R(R74) ,.T_L(T72), .T_R(T74), .R_old(R_old), .Z(Z73), .R(R73), .T(T73));
medianFilterCell  m74(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z73), .R_L(R73),.R_R(R75) ,.T_L(T73), .T_R(T75), .R_old(R_old), .Z(Z74), .R(R74), .T(T74));
medianFilterCell  m75(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z74), .R_L(R74),.R_R(R76) ,.T_L(T74), .T_R(T76), .R_old(R_old), .Z(Z75), .R(R75), .T(T75));
medianFilterCell  m76(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z75), .R_L(R75),.R_R(R77) ,.T_L(T75), .T_R(T77), .R_old(R_old), .Z(Z76), .R(R76), .T(T76));
medianFilterCell  m77(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z76), .R_L(R76),.R_R(R78) ,.T_L(T76), .T_R(T78), .R_old(R_old), .Z(Z77), .R(R77), .T(T77));
medianFilterCell  m78(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z77), .R_L(R77),.R_R(R79) ,.T_L(T77), .T_R(T79), .R_old(R_old), .Z(Z78), .R(R78), .T(T78));
medianFilterCell  m79(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z78), .R_L(R78),.R_R(R80) ,.T_L(T78), .T_R(T80), .R_old(R_old), .Z(Z79), .R(R79), .T(T79));
medianFilterCell  m80(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z79), .R_L(R79),.R_R(R81) ,.T_L(T79), .T_R(T81), .R_old(R_old), .Z(Z80), .R(R80), .T(T80));
medianFilterCell  m81(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z80), .R_L(R80),.R_R(R82) ,.T_L(T80), .T_R(T82), .R_old(R_old), .Z(Z81), .R(R81), .T(T81));
medianFilterCell  m82(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z81), .R_L(R81),.R_R(R83) ,.T_L(T81), .T_R(T83), .R_old(R_old), .Z(Z82), .R(R82), .T(T82));
medianFilterCell  m83(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z82), .R_L(R82),.R_R(R84) ,.T_L(T82), .T_R(T84), .R_old(R_old), .Z(Z83), .R(R83), .T(T83));
medianFilterCell  m84(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z83), .R_L(R83),.R_R(R85) ,.T_L(T83), .T_R(T85), .R_old(R_old), .Z(Z84), .R(R84), .T(T84));
medianFilterCell  m85(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z84), .R_L(R84),.R_R(R86) ,.T_L(T84), .T_R(T86), .R_old(R_old), .Z(Z85), .R(R85), .T(T85));
medianFilterCell  m86(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z85), .R_L(R85),.R_R(R87) ,.T_L(T85), .T_R(T87), .R_old(R_old), .Z(Z86), .R(R86), .T(T86));
medianFilterCell  m87(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z86), .R_L(R86),.R_R(R88) ,.T_L(T86), .T_R(T88), .R_old(R_old), .Z(Z87), .R(R87), .T(T87));
medianFilterCell  m88(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z87), .R_L(R87),.R_R(R89) ,.T_L(T87), .T_R(T89), .R_old(R_old), .Z(Z88), .R(R88), .T(T88));
medianFilterCell  m89(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z88), .R_L(R88),.R_R(R90) ,.T_L(T88), .T_R(T90), .R_old(R_old), .Z(Z89), .R(R89), .T(T89));
medianFilterCell  m90(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z89), .R_L(R89),.R_R(R91) ,.T_L(T89), .T_R(T91), .R_old(R_old), .Z(Z90), .R(R90), .T(T90));
medianFilterCell  m91(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z90), .R_L(R90),.R_R(R92) ,.T_L(T90), .T_R(T92), .R_old(R_old), .Z(Z91), .R(R91), .T(T91));
medianFilterCell  m92(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z91), .R_L(R91),.R_R(R93) ,.T_L(T91), .T_R(T93), .R_old(R_old), .Z(Z92), .R(R92), .T(T92));
medianFilterCell  m93(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z92), .R_L(R92),.R_R(R94) ,.T_L(T92), .T_R(T94), .R_old(R_old), .Z(Z93), .R(R93), .T(T93));
medianFilterCell  m94(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z93), .R_L(R93),.R_R(R95) ,.T_L(T93), .T_R(T95), .R_old(R_old), .Z(Z94), .R(R94), .T(T94));
medianFilterCell  m95(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z94), .R_L(R94),.R_R(R96) ,.T_L(T94), .T_R(T96), .R_old(R_old), .Z(Z95), .R(R95), .T(T95));
medianFilterCell  m96(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z95), .R_L(R95),.R_R(R97) ,.T_L(T95), .T_R(T97), .R_old(R_old), .Z(Z96), .R(R96), .T(T96));
medianFilterCell  m97(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z96), .R_L(R96),.R_R(R98) ,.T_L(T96), .T_R(T98), .R_old(R_old), .Z(Z97), .R(R97), .T(T97));
medianFilterCell  m98(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z97), .R_L(R97),.R_R(R99) ,.T_L(T97), .T_R(T99), .R_old(R_old), .Z(Z98), .R(R98), .T(T98));
medianFilterCell  m99(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z98), .R_L(R98),.R_R(R100) ,.T_L(T98), .T_R(T100), .R_old(R_old), .Z(Z99), .R(R99), .T(T99));
medianFilterCell  m100(.X(X) ,.clk(clk), .reset(reset) ,.Z_L(Z99), .R_L(R99),.R_R(R101) ,.T_L(T99), .T_R(T101), .R_old(R_old), .Z(Z100), .R(R100), .T(T100));
medianCell_rightMst  m101(.X(X) ,.clk(clk), .reset(reset), .Z_L(Z100), .R_L(R100), .T_L(T100), .R_old(R_old), .R(R101),.T(T101));


endmodule