`timescale 1ns / 1ps

module MatrixAdd_10_12_10PV_noHR_NIR_AXIStream
#(
parameter IN_DATA_LENGHT= 3840, 
parameter OUT_DATA_LENGHT= 2040 
)( 

input aclk,
input aresetn,
input enable,
input [IN_DATA_LENGHT-1:0]s_axi_data,
input s_axi_valid,
input m_axi_ready,
output reg[OUT_DATA_LENGHT-1:0]m_axi_data,
output reg m_axi_valid,
output reg s_axi_ready
);

reg inready;
reg [IN_DATA_LENGHT-1:0]indata;
wire outready;
wire earlyoutready;
wire [OUT_DATA_LENGHT-1:0]outdata;
////////////////instancing wrapping module///////////////////
MatrixAdd_10_12_10PV_noHR_NIR MatrixAdd_10_12_10PV_noHR_NIR_inst(
.clk(aclk),
.reset(!aresetn),
.enable(enable),
.inReady(inready),
.A0V0(indata[3839:3824]),
.A1V0(indata[3823:3808]),
.A2V0(indata[3807:3792]),
.A3V0(indata[3791:3776]),
.A4V0(indata[3775:3760]),
.A5V0(indata[3759:3744]),
.A6V0(indata[3743:3728]),
.A7V0(indata[3727:3712]),
.A8V0(indata[3711:3696]),
.A9V0(indata[3695:3680]),
.A10V0(indata[3679:3664]),
.A11V0(indata[3663:3648]),
.A0V1(indata[3647:3632]),
.A1V1(indata[3631:3616]),
.A2V1(indata[3615:3600]),
.A3V1(indata[3599:3584]),
.A4V1(indata[3583:3568]),
.A5V1(indata[3567:3552]),
.A6V1(indata[3551:3536]),
.A7V1(indata[3535:3520]),
.A8V1(indata[3519:3504]),
.A9V1(indata[3503:3488]),
.A10V1(indata[3487:3472]),
.A11V1(indata[3471:3456]),
.A0V2(indata[3455:3440]),
.A1V2(indata[3439:3424]),
.A2V2(indata[3423:3408]),
.A3V2(indata[3407:3392]),
.A4V2(indata[3391:3376]),
.A5V2(indata[3375:3360]),
.A6V2(indata[3359:3344]),
.A7V2(indata[3343:3328]),
.A8V2(indata[3327:3312]),
.A9V2(indata[3311:3296]),
.A10V2(indata[3295:3280]),
.A11V2(indata[3279:3264]),
.A0V3(indata[3263:3248]),
.A1V3(indata[3247:3232]),
.A2V3(indata[3231:3216]),
.A3V3(indata[3215:3200]),
.A4V3(indata[3199:3184]),
.A5V3(indata[3183:3168]),
.A6V3(indata[3167:3152]),
.A7V3(indata[3151:3136]),
.A8V3(indata[3135:3120]),
.A9V3(indata[3119:3104]),
.A10V3(indata[3103:3088]),
.A11V3(indata[3087:3072]),
.A0V4(indata[3071:3056]),
.A1V4(indata[3055:3040]),
.A2V4(indata[3039:3024]),
.A3V4(indata[3023:3008]),
.A4V4(indata[3007:2992]),
.A5V4(indata[2991:2976]),
.A6V4(indata[2975:2960]),
.A7V4(indata[2959:2944]),
.A8V4(indata[2943:2928]),
.A9V4(indata[2927:2912]),
.A10V4(indata[2911:2896]),
.A11V4(indata[2895:2880]),
.A0V5(indata[2879:2864]),
.A1V5(indata[2863:2848]),
.A2V5(indata[2847:2832]),
.A3V5(indata[2831:2816]),
.A4V5(indata[2815:2800]),
.A5V5(indata[2799:2784]),
.A6V5(indata[2783:2768]),
.A7V5(indata[2767:2752]),
.A8V5(indata[2751:2736]),
.A9V5(indata[2735:2720]),
.A10V5(indata[2719:2704]),
.A11V5(indata[2703:2688]),
.A0V6(indata[2687:2672]),
.A1V6(indata[2671:2656]),
.A2V6(indata[2655:2640]),
.A3V6(indata[2639:2624]),
.A4V6(indata[2623:2608]),
.A5V6(indata[2607:2592]),
.A6V6(indata[2591:2576]),
.A7V6(indata[2575:2560]),
.A8V6(indata[2559:2544]),
.A9V6(indata[2543:2528]),
.A10V6(indata[2527:2512]),
.A11V6(indata[2511:2496]),
.A0V7(indata[2495:2480]),
.A1V7(indata[2479:2464]),
.A2V7(indata[2463:2448]),
.A3V7(indata[2447:2432]),
.A4V7(indata[2431:2416]),
.A5V7(indata[2415:2400]),
.A6V7(indata[2399:2384]),
.A7V7(indata[2383:2368]),
.A8V7(indata[2367:2352]),
.A9V7(indata[2351:2336]),
.A10V7(indata[2335:2320]),
.A11V7(indata[2319:2304]),
.A0V8(indata[2303:2288]),
.A1V8(indata[2287:2272]),
.A2V8(indata[2271:2256]),
.A3V8(indata[2255:2240]),
.A4V8(indata[2239:2224]),
.A5V8(indata[2223:2208]),
.A6V8(indata[2207:2192]),
.A7V8(indata[2191:2176]),
.A8V8(indata[2175:2160]),
.A9V8(indata[2159:2144]),
.A10V8(indata[2143:2128]),
.A11V8(indata[2127:2112]),
.A0V9(indata[2111:2096]),
.A1V9(indata[2095:2080]),
.A2V9(indata[2079:2064]),
.A3V9(indata[2063:2048]),
.A4V9(indata[2047:2032]),
.A5V9(indata[2031:2016]),
.A6V9(indata[2015:2000]),
.A7V9(indata[1999:1984]),
.A8V9(indata[1983:1968]),
.A9V9(indata[1967:1952]),
.A10V9(indata[1951:1936]),
.A11V9(indata[1935:1920]),
.B0V0(indata[1919:1904]),
.B1V0(indata[1903:1888]),
.B2V0(indata[1887:1872]),
.B3V0(indata[1871:1856]),
.B4V0(indata[1855:1840]),
.B5V0(indata[1839:1824]),
.B6V0(indata[1823:1808]),
.B7V0(indata[1807:1792]),
.B8V0(indata[1791:1776]),
.B9V0(indata[1775:1760]),
.B10V0(indata[1759:1744]),
.B11V0(indata[1743:1728]),
.B0V1(indata[1727:1712]),
.B1V1(indata[1711:1696]),
.B2V1(indata[1695:1680]),
.B3V1(indata[1679:1664]),
.B4V1(indata[1663:1648]),
.B5V1(indata[1647:1632]),
.B6V1(indata[1631:1616]),
.B7V1(indata[1615:1600]),
.B8V1(indata[1599:1584]),
.B9V1(indata[1583:1568]),
.B10V1(indata[1567:1552]),
.B11V1(indata[1551:1536]),
.B0V2(indata[1535:1520]),
.B1V2(indata[1519:1504]),
.B2V2(indata[1503:1488]),
.B3V2(indata[1487:1472]),
.B4V2(indata[1471:1456]),
.B5V2(indata[1455:1440]),
.B6V2(indata[1439:1424]),
.B7V2(indata[1423:1408]),
.B8V2(indata[1407:1392]),
.B9V2(indata[1391:1376]),
.B10V2(indata[1375:1360]),
.B11V2(indata[1359:1344]),
.B0V3(indata[1343:1328]),
.B1V3(indata[1327:1312]),
.B2V3(indata[1311:1296]),
.B3V3(indata[1295:1280]),
.B4V3(indata[1279:1264]),
.B5V3(indata[1263:1248]),
.B6V3(indata[1247:1232]),
.B7V3(indata[1231:1216]),
.B8V3(indata[1215:1200]),
.B9V3(indata[1199:1184]),
.B10V3(indata[1183:1168]),
.B11V3(indata[1167:1152]),
.B0V4(indata[1151:1136]),
.B1V4(indata[1135:1120]),
.B2V4(indata[1119:1104]),
.B3V4(indata[1103:1088]),
.B4V4(indata[1087:1072]),
.B5V4(indata[1071:1056]),
.B6V4(indata[1055:1040]),
.B7V4(indata[1039:1024]),
.B8V4(indata[1023:1008]),
.B9V4(indata[1007:992]),
.B10V4(indata[991:976]),
.B11V4(indata[975:960]),
.B0V5(indata[959:944]),
.B1V5(indata[943:928]),
.B2V5(indata[927:912]),
.B3V5(indata[911:896]),
.B4V5(indata[895:880]),
.B5V5(indata[879:864]),
.B6V5(indata[863:848]),
.B7V5(indata[847:832]),
.B8V5(indata[831:816]),
.B9V5(indata[815:800]),
.B10V5(indata[799:784]),
.B11V5(indata[783:768]),
.B0V6(indata[767:752]),
.B1V6(indata[751:736]),
.B2V6(indata[735:720]),
.B3V6(indata[719:704]),
.B4V6(indata[703:688]),
.B5V6(indata[687:672]),
.B6V6(indata[671:656]),
.B7V6(indata[655:640]),
.B8V6(indata[639:624]),
.B9V6(indata[623:608]),
.B10V6(indata[607:592]),
.B11V6(indata[591:576]),
.B0V7(indata[575:560]),
.B1V7(indata[559:544]),
.B2V7(indata[543:528]),
.B3V7(indata[527:512]),
.B4V7(indata[511:496]),
.B5V7(indata[495:480]),
.B6V7(indata[479:464]),
.B7V7(indata[463:448]),
.B8V7(indata[447:432]),
.B9V7(indata[431:416]),
.B10V7(indata[415:400]),
.B11V7(indata[399:384]),
.B0V8(indata[383:368]),
.B1V8(indata[367:352]),
.B2V8(indata[351:336]),
.B3V8(indata[335:320]),
.B4V8(indata[319:304]),
.B5V8(indata[303:288]),
.B6V8(indata[287:272]),
.B7V8(indata[271:256]),
.B8V8(indata[255:240]),
.B9V8(indata[239:224]),
.B10V8(indata[223:208]),
.B11V8(indata[207:192]),
.B0V9(indata[191:176]),
.B1V9(indata[175:160]),
.B2V9(indata[159:144]),
.B3V9(indata[143:128]),
.B4V9(indata[127:112]),
.B5V9(indata[111:96]),
.B6V9(indata[95:80]),
.B7V9(indata[79:64]),
.B8V9(indata[63:48]),
.B9V9(indata[47:32]),
.B10V9(indata[31:16]),
.B11V9(indata[15:0]),
.V0toV11outReady(outready),
.S0V0(outdata[2039:2024]),
.S1V0(outdata[2023:2008]),
.S2V0(outdata[2007:1992]),
.S3V0(outdata[1991:1976]),
.S4V0(outdata[1975:1960]),
.S5V0(outdata[1959:1944]),
.S6V0(outdata[1943:1928]),
.S7V0(outdata[1927:1912]),
.S8V0(outdata[1911:1896]),
.S9V0(outdata[1895:1880]),
.S10V0(outdata[1879:1864]),
.S11V0(outdata[1863:1848]),
.S0V1(outdata[1847:1832]),
.S1V1(outdata[1831:1816]),
.S2V1(outdata[1815:1800]),
.S3V1(outdata[1799:1784]),
.S4V1(outdata[1783:1768]),
.S5V1(outdata[1767:1752]),
.S6V1(outdata[1751:1736]),
.S7V1(outdata[1735:1720]),
.S8V1(outdata[1719:1704]),
.S9V1(outdata[1703:1688]),
.S10V1(outdata[1687:1672]),
.S11V1(outdata[1671:1656]),
.S0V2(outdata[1655:1640]),
.S1V2(outdata[1639:1624]),
.S2V2(outdata[1623:1608]),
.S3V2(outdata[1607:1592]),
.S4V2(outdata[1591:1576]),
.S5V2(outdata[1575:1560]),
.S6V2(outdata[1559:1544]),
.S7V2(outdata[1543:1528]),
.S8V2(outdata[1527:1512]),
.S9V2(outdata[1511:1496]),
.S10V2(outdata[1495:1480]),
.S11V2(outdata[1479:1464]),
.S0V3(outdata[1463:1448]),
.S1V3(outdata[1447:1432]),
.S2V3(outdata[1431:1416]),
.S3V3(outdata[1415:1400]),
.S4V3(outdata[1399:1384]),
.S5V3(outdata[1383:1368]),
.S6V3(outdata[1367:1352]),
.S7V3(outdata[1351:1336]),
.S8V3(outdata[1335:1320]),
.S9V3(outdata[1319:1304]),
.S10V3(outdata[1303:1288]),
.S11V3(outdata[1287:1272]),
.S0V4(outdata[1271:1256]),
.S1V4(outdata[1255:1240]),
.S2V4(outdata[1239:1224]),
.S3V4(outdata[1223:1208]),
.S4V4(outdata[1207:1192]),
.S5V4(outdata[1191:1176]),
.S6V4(outdata[1175:1160]),
.S7V4(outdata[1159:1144]),
.S8V4(outdata[1143:1128]),
.S9V4(outdata[1127:1112]),
.S10V4(outdata[1111:1096]),
.S11V4(outdata[1095:1080]),
.S0V5(outdata[1079:1064]),
.S1V5(outdata[1063:1048]),
.S2V5(outdata[1047:1032]),
.S3V5(outdata[1031:1016]),
.S4V5(outdata[1015:1000]),
.S5V5(outdata[999:984]),
.S6V5(outdata[983:968]),
.S7V5(outdata[967:952]),
.S8V5(outdata[951:936]),
.S9V5(outdata[935:920]),
.S10V5(outdata[919:904]),
.S11V5(outdata[903:888]),
.S0V6(outdata[887:872]),
.S1V6(outdata[871:856]),
.S2V6(outdata[855:840]),
.S3V6(outdata[839:824]),
.S4V6(outdata[823:808]),
.S5V6(outdata[807:792]),
.S6V6(outdata[791:776]),
.S7V6(outdata[775:760]),
.S8V6(outdata[759:744]),
.S9V6(outdata[743:728]),
.S10V6(outdata[727:712]),
.S11V6(outdata[711:696]),
.S0V7(outdata[695:680]),
.S1V7(outdata[679:664]),
.S2V7(outdata[663:648]),
.S3V7(outdata[647:632]),
.S4V7(outdata[631:616]),
.S5V7(outdata[615:600]),
.S6V7(outdata[599:584]),
.S7V7(outdata[583:568]),
.S8V7(outdata[567:552]),
.S9V7(outdata[551:536]),
.S10V7(outdata[535:520]),
.S11V7(outdata[519:504]),
.S0V8(outdata[503:488]),
.S1V8(outdata[487:472]),
.S2V8(outdata[471:456]),
.S3V8(outdata[455:440]),
.S4V8(outdata[439:424]),
.S5V8(outdata[423:408]),
.S6V8(outdata[407:392]),
.S7V8(outdata[391:376]),
.S8V8(outdata[375:360]),
.S9V8(outdata[359:344]),
.S10V8(outdata[343:328]),
.S11V8(outdata[327:312]),
.S0V9(outdata[311:296]),
.S1V9(outdata[295:280]),
.S2V9(outdata[279:264]),
.S3V9(outdata[263:248]),
.S4V9(outdata[247:232]),
.S5V9(outdata[231:216]),
.S6V9(outdata[215:200]),
.S7V9(outdata[199:184]),
.S8V9(outdata[183:168]),
.S9V9(outdata[167:152]),
.S10V9(outdata[151:136]),
.S11V9(outdata[135:120]),
.V0toV12earlyOutReady(earlyoutready)
);
/////////////////Main body/////////////
always @(posedge aclk)begin
 if(aresetn==0)begin
  m_axi_data<=0;
  m_axi_valid<=0;
 end
 else begin
  if(m_axi_ready==1 && m_axi_valid==1)begin
   m_axi_valid<=0;
  end
  else if(outready==1)begin
   m_axi_valid<=1;
   m_axi_data<=outdata;
  end
 end
end
always @(posedge aclk)begin
 if(aresetn==0)begin
  s_axi_ready<=1;
  inready<=0;
  indata<=0;
 end
 else begin
  inready<=0;
  if(s_axi_valid==1 && s_axi_ready==1)begin
   s_axi_ready<=0;
   inready<=1;
   indata<= s_axi_data;
  end
  else if(m_axi_valid==1 && m_axi_ready==1)begin
   s_axi_ready<=1;
  end
 end
end

endmodule
