`timescale 1ns / 1ps

module MatrixAdd_12_10_12PV_noHR_NIR
#(
parameter IN_WIDTH = 16
)(
input clk, reset, enable,
output reg vectorSetInNo = 0,
input inReady,
input signed [IN_WIDTH-1:0] A0V0, A1V0, A2V0, A3V0, A4V0, A5V0, A6V0, A7V0, A8V0, A9V0, 
A0V1, A1V1, A2V1, A3V1, A4V1, A5V1, A6V1, A7V1, A8V1, A9V1, 
A0V2, A1V2, A2V2, A3V2, A4V2, A5V2, A6V2, A7V2, A8V2, A9V2, 
A0V3, A1V3, A2V3, A3V3, A4V3, A5V3, A6V3, A7V3, A8V3, A9V3, 
A0V4, A1V4, A2V4, A3V4, A4V4, A5V4, A6V4, A7V4, A8V4, A9V4, 
A0V5, A1V5, A2V5, A3V5, A4V5, A5V5, A6V5, A7V5, A8V5, A9V5, 
A0V6, A1V6, A2V6, A3V6, A4V6, A5V6, A6V6, A7V6, A8V6, A9V6, 
A0V7, A1V7, A2V7, A3V7, A4V7, A5V7, A6V7, A7V7, A8V7, A9V7, 
A0V8, A1V8, A2V8, A3V8, A4V8, A5V8, A6V8, A7V8, A8V8, A9V8, 
A0V9, A1V9, A2V9, A3V9, A4V9, A5V9, A6V9, A7V9, A8V9, A9V9, 
A0V10, A1V10, A2V10, A3V10, A4V10, A5V10, A6V10, A7V10, A8V10, A9V10, 
A0V11, A1V11, A2V11, A3V11, A4V11, A5V11, A6V11, A7V11, A8V11, A9V11, 
input signed [IN_WIDTH-1:0] B0V0, B1V0, B2V0, B3V0, B4V0, B5V0, B6V0, B7V0, B8V0, B9V0, 
B0V1, B1V1, B2V1, B3V1, B4V1, B5V1, B6V1, B7V1, B8V1, B9V1, 
B0V2, B1V2, B2V2, B3V2, B4V2, B5V2, B6V2, B7V2, B8V2, B9V2, 
B0V3, B1V3, B2V3, B3V3, B4V3, B5V3, B6V3, B7V3, B8V3, B9V3, 
B0V4, B1V4, B2V4, B3V4, B4V4, B5V4, B6V4, B7V4, B8V4, B9V4, 
B0V5, B1V5, B2V5, B3V5, B4V5, B5V5, B6V5, B7V5, B8V5, B9V5, 
B0V6, B1V6, B2V6, B3V6, B4V6, B5V6, B6V6, B7V6, B8V6, B9V6, 
B0V7, B1V7, B2V7, B3V7, B4V7, B5V7, B6V7, B7V7, B8V7, B9V7, 
B0V8, B1V8, B2V8, B3V8, B4V8, B5V8, B6V8, B7V8, B8V8, B9V8, 
B0V9, B1V9, B2V9, B3V9, B4V9, B5V9, B6V9, B7V9, B8V9, B9V9, 
B0V10, B1V10, B2V10, B3V10, B4V10, B5V10, B6V10, B7V10, B8V10, B9V10, 
B0V11, B1V11, B2V11, B3V11, B4V11, B5V11, B6V11, B7V11, B8V11, B9V11, 
output V0toV11outReady,
output reg VNoutReady1 = 0, //not used
output reg VNoutReady2 = 0, //not used
output reg vectorSetOutNo = 1,
output signed [IN_WIDTH:0] S0V0, S1V0, S2V0, S3V0, S4V0, S5V0, S6V0, S7V0, S8V0, S9V0, 
S0V1, S1V1, S2V1, S3V1, S4V1, S5V1, S6V1, S7V1, S8V1, S9V1, 
S0V2, S1V2, S2V2, S3V2, S4V2, S5V2, S6V2, S7V2, S8V2, S9V2, 
S0V3, S1V3, S2V3, S3V3, S4V3, S5V3, S6V3, S7V3, S8V3, S9V3, 
S0V4, S1V4, S2V4, S3V4, S4V4, S5V4, S6V4, S7V4, S8V4, S9V4, 
S0V5, S1V5, S2V5, S3V5, S4V5, S5V5, S6V5, S7V5, S8V5, S9V5, 
S0V6, S1V6, S2V6, S3V6, S4V6, S5V6, S6V6, S7V6, S8V6, S9V6, 
S0V7, S1V7, S2V7, S3V7, S4V7, S5V7, S6V7, S7V7, S8V7, S9V7, 
S0V8, S1V8, S2V8, S3V8, S4V8, S5V8, S6V8, S7V8, S8V8, S9V8, 
S0V9, S1V9, S2V9, S3V9, S4V9, S5V9, S6V9, S7V9, S8V9, S9V9, 
S0V10, S1V10, S2V10, S3V10, S4V10, S5V10, S6V10, S7V10, S8V10, S9V10, 
S0V11, S1V11, S2V11, S3V11, S4V11, S5V11, S6V11, S7V11, S8V11, S9V11, 
output V0toV11earlyOutReady,
output reg CNearlyOutReady1 = 0, //not used
output reg CNearlyOutReady2 = 0 //not used
);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_0(clk, reset, enable,
	inReady,
	A0V0, A1V0, A2V0, A3V0, A4V0, A5V0, A6V0, A7V0, A8V0, A9V0, 
	B0V0, B1V0, B2V0, B3V0, B4V0, B5V0, B6V0, B7V0, B8V0, B9V0, 
	V0toV11outReady,
	S0V0, S1V0, S2V0, S3V0, S4V0, S5V0, S6V0, S7V0, S8V0, S9V0, 
	V0toV11earlyOutReady
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_1(clk, reset, enable,
	inReady,
	A0V1, A1V1, A2V1, A3V1, A4V1, A5V1, A6V1, A7V1, A8V1, A9V1, 
	B0V1, B1V1, B2V1, B3V1, B4V1, B5V1, B6V1, B7V1, B8V1, B9V1, 
	VA1OR, //not used
	S0V1, S1V1, S2V1, S3V1, S4V1, S5V1, S6V1, S7V1, S8V1, S9V1, 
	VA1EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_2(clk, reset, enable,
	inReady,
	A0V2, A1V2, A2V2, A3V2, A4V2, A5V2, A6V2, A7V2, A8V2, A9V2, 
	B0V2, B1V2, B2V2, B3V2, B4V2, B5V2, B6V2, B7V2, B8V2, B9V2, 
	VA2OR, //not used
	S0V2, S1V2, S2V2, S3V2, S4V2, S5V2, S6V2, S7V2, S8V2, S9V2, 
	VA2EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_3(clk, reset, enable,
	inReady,
	A0V3, A1V3, A2V3, A3V3, A4V3, A5V3, A6V3, A7V3, A8V3, A9V3, 
	B0V3, B1V3, B2V3, B3V3, B4V3, B5V3, B6V3, B7V3, B8V3, B9V3, 
	VA3OR, //not used
	S0V3, S1V3, S2V3, S3V3, S4V3, S5V3, S6V3, S7V3, S8V3, S9V3, 
	VA3EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_4(clk, reset, enable,
	inReady,
	A0V4, A1V4, A2V4, A3V4, A4V4, A5V4, A6V4, A7V4, A8V4, A9V4, 
	B0V4, B1V4, B2V4, B3V4, B4V4, B5V4, B6V4, B7V4, B8V4, B9V4, 
	VA4OR, //not used
	S0V4, S1V4, S2V4, S3V4, S4V4, S5V4, S6V4, S7V4, S8V4, S9V4, 
	VA4EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_5(clk, reset, enable,
	inReady,
	A0V5, A1V5, A2V5, A3V5, A4V5, A5V5, A6V5, A7V5, A8V5, A9V5, 
	B0V5, B1V5, B2V5, B3V5, B4V5, B5V5, B6V5, B7V5, B8V5, B9V5, 
	VA5OR, //not used
	S0V5, S1V5, S2V5, S3V5, S4V5, S5V5, S6V5, S7V5, S8V5, S9V5, 
	VA5EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_6(clk, reset, enable,
	inReady,
	A0V6, A1V6, A2V6, A3V6, A4V6, A5V6, A6V6, A7V6, A8V6, A9V6, 
	B0V6, B1V6, B2V6, B3V6, B4V6, B5V6, B6V6, B7V6, B8V6, B9V6, 
	VA6OR, //not used
	S0V6, S1V6, S2V6, S3V6, S4V6, S5V6, S6V6, S7V6, S8V6, S9V6, 
	VA6EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_7(clk, reset, enable,
	inReady,
	A0V7, A1V7, A2V7, A3V7, A4V7, A5V7, A6V7, A7V7, A8V7, A9V7, 
	B0V7, B1V7, B2V7, B3V7, B4V7, B5V7, B6V7, B7V7, B8V7, B9V7, 
	VA7OR, //not used
	S0V7, S1V7, S2V7, S3V7, S4V7, S5V7, S6V7, S7V7, S8V7, S9V7, 
	VA7EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_8(clk, reset, enable,
	inReady,
	A0V8, A1V8, A2V8, A3V8, A4V8, A5V8, A6V8, A7V8, A8V8, A9V8, 
	B0V8, B1V8, B2V8, B3V8, B4V8, B5V8, B6V8, B7V8, B8V8, B9V8, 
	VA8OR, //not used
	S0V8, S1V8, S2V8, S3V8, S4V8, S5V8, S6V8, S7V8, S8V8, S9V8, 
	VA8EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_9(clk, reset, enable,
	inReady,
	A0V9, A1V9, A2V9, A3V9, A4V9, A5V9, A6V9, A7V9, A8V9, A9V9, 
	B0V9, B1V9, B2V9, B3V9, B4V9, B5V9, B6V9, B7V9, B8V9, B9V9, 
	VA9OR, //not used
	S0V9, S1V9, S2V9, S3V9, S4V9, S5V9, S6V9, S7V9, S8V9, S9V9, 
	VA9EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_10(clk, reset, enable,
	inReady,
	A0V10, A1V10, A2V10, A3V10, A4V10, A5V10, A6V10, A7V10, A8V10, A9V10, 
	B0V10, B1V10, B2V10, B3V10, B4V10, B5V10, B6V10, B7V10, B8V10, B9V10, 
	VA10OR, //not used
	S0V10, S1V10, S2V10, S3V10, S4V10, S5V10, S6V10, S7V10, S8V10, S9V10, 
	VA10EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_11(clk, reset, enable,
	inReady,
	A0V11, A1V11, A2V11, A3V11, A4V11, A5V11, A6V11, A7V11, A8V11, A9V11, 
	B0V11, B1V11, B2V11, B3V11, B4V11, B5V11, B6V11, B7V11, B8V11, B9V11, 
	VA11OR, //not used
	S0V11, S1V11, S2V11, S3V11, S4V11, S5V11, S6V11, S7V11, S8V11, S9V11, 
	VA11EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_0(clk, reset, enable,
	inReady,
	A0V0, A1V0, A2V0, A3V0, A4V0, A5V0, A6V0, A7V0, A8V0, A9V0, 
	B0V0, B1V0, B2V0, B3V0, B4V0, B5V0, B6V0, B7V0, B8V0, B9V0, 
	V0toV11outReady,
	S0V0, S1V0, S2V0, S3V0, S4V0, S5V0, S6V0, S7V0, S8V0, S9V0, 
	V0toV11earlyOutReady
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_1(clk, reset, enable,
	inReady,
	A0V1, A1V1, A2V1, A3V1, A4V1, A5V1, A6V1, A7V1, A8V1, A9V1, 
	B0V1, B1V1, B2V1, B3V1, B4V1, B5V1, B6V1, B7V1, B8V1, B9V1, 
	VA1OR, //not used
	S0V1, S1V1, S2V1, S3V1, S4V1, S5V1, S6V1, S7V1, S8V1, S9V1, 
	VA1EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_2(clk, reset, enable,
	inReady,
	A0V2, A1V2, A2V2, A3V2, A4V2, A5V2, A6V2, A7V2, A8V2, A9V2, 
	B0V2, B1V2, B2V2, B3V2, B4V2, B5V2, B6V2, B7V2, B8V2, B9V2, 
	VA2OR, //not used
	S0V2, S1V2, S2V2, S3V2, S4V2, S5V2, S6V2, S7V2, S8V2, S9V2, 
	VA2EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_3(clk, reset, enable,
	inReady,
	A0V3, A1V3, A2V3, A3V3, A4V3, A5V3, A6V3, A7V3, A8V3, A9V3, 
	B0V3, B1V3, B2V3, B3V3, B4V3, B5V3, B6V3, B7V3, B8V3, B9V3, 
	VA3OR, //not used
	S0V3, S1V3, S2V3, S3V3, S4V3, S5V3, S6V3, S7V3, S8V3, S9V3, 
	VA3EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_4(clk, reset, enable,
	inReady,
	A0V4, A1V4, A2V4, A3V4, A4V4, A5V4, A6V4, A7V4, A8V4, A9V4, 
	B0V4, B1V4, B2V4, B3V4, B4V4, B5V4, B6V4, B7V4, B8V4, B9V4, 
	VA4OR, //not used
	S0V4, S1V4, S2V4, S3V4, S4V4, S5V4, S6V4, S7V4, S8V4, S9V4, 
	VA4EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_5(clk, reset, enable,
	inReady,
	A0V5, A1V5, A2V5, A3V5, A4V5, A5V5, A6V5, A7V5, A8V5, A9V5, 
	B0V5, B1V5, B2V5, B3V5, B4V5, B5V5, B6V5, B7V5, B8V5, B9V5, 
	VA5OR, //not used
	S0V5, S1V5, S2V5, S3V5, S4V5, S5V5, S6V5, S7V5, S8V5, S9V5, 
	VA5EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_6(clk, reset, enable,
	inReady,
	A0V6, A1V6, A2V6, A3V6, A4V6, A5V6, A6V6, A7V6, A8V6, A9V6, 
	B0V6, B1V6, B2V6, B3V6, B4V6, B5V6, B6V6, B7V6, B8V6, B9V6, 
	VA6OR, //not used
	S0V6, S1V6, S2V6, S3V6, S4V6, S5V6, S6V6, S7V6, S8V6, S9V6, 
	VA6EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_7(clk, reset, enable,
	inReady,
	A0V7, A1V7, A2V7, A3V7, A4V7, A5V7, A6V7, A7V7, A8V7, A9V7, 
	B0V7, B1V7, B2V7, B3V7, B4V7, B5V7, B6V7, B7V7, B8V7, B9V7, 
	VA7OR, //not used
	S0V7, S1V7, S2V7, S3V7, S4V7, S5V7, S6V7, S7V7, S8V7, S9V7, 
	VA7EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_8(clk, reset, enable,
	inReady,
	A0V8, A1V8, A2V8, A3V8, A4V8, A5V8, A6V8, A7V8, A8V8, A9V8, 
	B0V8, B1V8, B2V8, B3V8, B4V8, B5V8, B6V8, B7V8, B8V8, B9V8, 
	VA8OR, //not used
	S0V8, S1V8, S2V8, S3V8, S4V8, S5V8, S6V8, S7V8, S8V8, S9V8, 
	VA8EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_9(clk, reset, enable,
	inReady,
	A0V9, A1V9, A2V9, A3V9, A4V9, A5V9, A6V9, A7V9, A8V9, A9V9, 
	B0V9, B1V9, B2V9, B3V9, B4V9, B5V9, B6V9, B7V9, B8V9, B9V9, 
	VA9OR, //not used
	S0V9, S1V9, S2V9, S3V9, S4V9, S5V9, S6V9, S7V9, S8V9, S9V9, 
	VA9EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_10(clk, reset, enable,
	inReady,
	A0V10, A1V10, A2V10, A3V10, A4V10, A5V10, A6V10, A7V10, A8V10, A9V10, 
	B0V10, B1V10, B2V10, B3V10, B4V10, B5V10, B6V10, B7V10, B8V10, B9V10, 
	VA10OR, //not used
	S0V10, S1V10, S2V10, S3V10, S4V10, S5V10, S6V10, S7V10, S8V10, S9V10, 
	VA10EOR //not used
	);

VectorAdd_10_noHR_NIR#( .IN_WIDTH(IN_WIDTH) )
	VA_11(clk, reset, enable,
	inReady,
	A0V11, A1V11, A2V11, A3V11, A4V11, A5V11, A6V11, A7V11, A8V11, A9V11, 
	B0V11, B1V11, B2V11, B3V11, B4V11, B5V11, B6V11, B7V11, B8V11, B9V11, 
	VA11OR, //not used
	S0V11, S1V11, S2V11, S3V11, S4V11, S5V11, S6V11, S7V11, S8V11, S9V11, 
	VA11EOR //not used
	);

endmodule
