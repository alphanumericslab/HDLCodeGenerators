`timescale 1ns / 1ps
`include "macro.vh"
///////////////////////
module top ( clk ,reset ,X , W, median );

output [`DATA_LENGTH-1:0] median ;
input [`DATA_LENGTH-1:0] X;
input [`LOG_WMAX-1:0] W;
input clk ,reset ;

wire 	[`DATA_LENGTH-1:0] R_old ,R1_1 ,R2_1 ,R1_2 ,R2_2 ,R1_3 ,R2_3 ,R1_4 ,R2_4 ,R1_5 ,R2_5 ,R1_6 ,R2_6 ,R1_7 ,R2_7 ,R1_8 ,R2_8 ,R1_9 ,R2_9 ,R1_10 ,R2_10 ,R1_11 ,R2_11 ,R1_12 ,R2_12 ,R1_13 ,R2_13 ,R1_14 ,R2_14 ,R1_15 ,R2_15 ,R1_16 ,R2_16 ,R1_17 ,R2_17 ,R1_18 ,R2_18 ,R1_19 ,R2_19 ,R1_20 ,R2_20 ,R1_21 ,R2_21 ,R1_22 ,R2_22 ,R1_23 ,R2_23 ,R1_24 ,R2_24 ,R1_25 ,R2_25 ,R1_26 ,R2_26 ,R1_27 ,R2_27 ,R1_28 ,R2_28 ,R1_29 ,R2_29 ,R1_30 ,R2_30 ,R1_31 ,R2_31 ,R1_32 ,R2_32 ,R1_33 ,R2_33 ,R1_34 ,R2_34 ,R1_35 ,R2_35 ,R1_36 ,R2_36 ,R1_37 ,R2_37 ,R1_38 ,R2_38 ,R1_39 ,R2_39 ,R1_40 ,R2_40 ,R1_41 ,R2_41 ,R1_42 ,R2_42 ,R1_43 ,R2_43 ,R1_44 ,R2_44 ,R1_45 ,R2_45 ,R1_46 ,R2_46 ,R1_47 ,R2_47 ,R1_48 ,R2_48 ,R1_49 ,R2_49 ,R1_50 ,R2_50 ,R1_51 ,R2_51 ,R1_52 ,R2_52 ,R1_53 ,R2_53 ,R1_54 ,R2_54 ,R1_55 ,R2_55 ,R1_56 ,R2_56 ,R1_57 ,R2_57 ,R1_58 ,R2_58 ,R1_59 ,R2_59 ,R1_60 ,R2_60 ,R1_61 ,R2_61 ,R1_62 ,R2_62 ,R1_63 ,R2_63 ,R1_64 ,R2_64 ,R1_65 ,R2_65 ,R1_66 ,R2_66 ,R1_67 ,R2_67 ,R1_68 ,R2_68 ,R1_69 ,R2_69 ,R1_70 ,R2_70 ,R1_71 ,R2_71 ,R1_72 ,R2_72 ,R1_73 ,R2_73 ,R1_74 ,R2_74 ,R1_75 ,R2_75 ,R1_76 ,R2_76 ,R1_77 ,R2_77 ,R1_78 ,R2_78 ,R1_79 ,R2_79 ,R1_80 ,R2_80 ,R1_81 ,R2_81 ,R1_82 ,R2_82 ,R1_83 ,R2_83 ,R1_84 ,R2_84 ,R1_85 ,R2_85 ,R1_86 ,R2_86 ,R1_87 ,R2_87 ,R1_88 ,R2_88 ,R1_89 ,R2_89 ,R1_90 ,R2_90 ,R1_91 ,R2_91 ,R1_92 ,R2_92 ,R1_93 ,R2_93 ,R1_94 ,R2_94 ,R1_95 ,R2_95 ,R1_96 ,R2_96 ,R1_97 ,R2_97 ,R1_98 ,R2_98 ,R1_99 ,R2_99 ,R1_100 ,R2_100 ,R1_101 ,R2_101 ,R1_102 ,R2_102 ,R1_103 ,R2_103 ,R1_104 ,R2_104 ,R1_105 ,R2_105 ,R1_106 ,R2_106 ,R1_107 ,R2_107 ,R1_108 ,R2_108 ,R1_109 ,R2_109 ,R1_110 ,R2_110 ,R1_111 ,R2_111 ,R1_112 ,R2_112 ,R1_113 ,R2_113 ,R1_114 ,R2_114 ,R1_115 ,R2_115 ,R1_116 ,R2_116 ,R1_117 ,R2_117 ,R1_118 ,R2_118 ,R1_119 ,R2_119 ,R1_120 ,R2_120 ,R1_121 ,R2_121 ,R1_122 ,R2_122 ,R1_123 ,R2_123 ,R1_124 ,R2_124 ,R1_125 ,R2_125 ,R1_126 ,R2_126 ,R1_127 ,R2_127 ,R1_128 ,R2_128 ,R1_129 ,R2_129 ,R1_130 ,R2_130 ,R1_131 ,R2_131 ,R1_132 ,R2_132 ,R1_133 ,R2_133 ,R1_134 ,R2_134 ,R1_135 ,R2_135 ,R1_136 ,R2_136 ,R1_137 ,R2_137 ,R1_138 ,R2_138 ,R1_139 ,R2_139 ,R1_140 ,R2_140 ,R1_141 ,R2_141 ,R1_142 ,R2_142 ,R1_143 ,R2_143 ,R1_144 ,R2_144 ,R1_145 ,R2_145 ,R1_146 ,R2_146 ,R1_147 ,R2_147 ,R1_148 ,R2_148 ,R1_149 ,R2_149 ,R1_150 ,R2_150 ,R1_151 ,R2_151 ,R1_152 ,R2_152 ,R1_153 ,R2_153 ,R1_154 ,R2_154 ,R1_155 ,R2_155 ,R1_156 ,R2_156 ,R1_157 ,R2_157 ,R1_158 ,R2_158 ,R1_159 ,R2_159 ,R1_160 ,R2_160 ,R1_161 ,R2_161 ,R1_162 ,R2_162 ,R1_163 ,R2_163 ,R1_164 ,R2_164 ,R1_165 ,R2_165 ,R1_166 ,R2_166 ,R1_167 ,R2_167 ,R1_168 ,R2_168 ,R1_169 ,R2_169 ,R1_170 ,R2_170 ,R1_171 ,R2_171 ,R1_172 ,R2_172 ,R1_173 ,R2_173 ,R1_174 ,R2_174 ,R1_175 ,R2_175 ,R1_176 ,R2_176 ,R1_177 ,R2_177 ,R1_178 ,R2_178 ,R1_179 ,R2_179 ,R1_180 ,R2_180 ,R1_181 ,R2_181 ,R1_182 ,R2_182 ,R1_183 ,R2_183 ,R1_184 ,R2_184 ,R1_185 ,R2_185 ,R1_186 ,R2_186 ,R1_187 ,R2_187 ,R1_188 ,R2_188 ,R1_189 ,R2_189 ,R1_190 ,R2_190 ,R1_191 ,R2_191 ,R1_192 ,R2_192 ,R1_193 ,R2_193 ,R1_194 ,R2_194 ,R1_195 ,R2_195 ,R1_196 ,R2_196 ,R1_197 ,R2_197 ,R1_198 ,R2_198 ,R1_199 ,R2_199 ,R1_200 ,R2_200 ,R1_201 ,R2_201;
wire 	T1 ,T2 ,T3 ,T4 ,T5 ,T6 ,T7 ,T8 ,T9 ,T10 ,T11 ,T12 ,T13 ,T14 ,T15 ,T16 ,T17 ,T18 ,T19 ,T20 ,T21 ,T22 ,T23 ,T24 ,T25 ,T26 ,T27 ,T28 ,T29 ,T30 ,T31 ,T32 ,T33 ,T34 ,T35 ,T36 ,T37 ,T38 ,T39 ,T40 ,T41 ,T42 ,T43 ,T44 ,T45 ,T46 ,T47 ,T48 ,T49 ,T50 ,T51 ,T52 ,T53 ,T54 ,T55 ,T56 ,T57 ,T58 ,T59 ,T60 ,T61 ,T62 ,T63 ,T64 ,T65 ,T66 ,T67 ,T68 ,T69 ,T70 ,T71 ,T72 ,T73 ,T74 ,T75 ,T76 ,T77 ,T78 ,T79 ,T80 ,T81 ,T82 ,T83 ,T84 ,T85 ,T86 ,T87 ,T88 ,T89 ,T90 ,T91 ,T92 ,T93 ,T94 ,T95 ,T96 ,T97 ,T98 ,T99 ,T100 ,T101 ,T102 ,T103 ,T104 ,T105 ,T106 ,T107 ,T108 ,T109 ,T110 ,T111 ,T112 ,T113 ,T114 ,T115 ,T116 ,T117 ,T118 ,T119 ,T120 ,T121 ,T122 ,T123 ,T124 ,T125 ,T126 ,T127 ,T128 ,T129 ,T130 ,T131 ,T132 ,T133 ,T134 ,T135 ,T136 ,T137 ,T138 ,T139 ,T140 ,T141 ,T142 ,T143 ,T144 ,T145 ,T146 ,T147 ,T148 ,T149 ,T150 ,T151 ,T152 ,T153 ,T154 ,T155 ,T156 ,T157 ,T158 ,T159 ,T160 ,T161 ,T162 ,T163 ,T164 ,T165 ,T166 ,T167 ,T168 ,T169 ,T170 ,T171 ,T172 ,T173 ,T174 ,T175 ,T176 ,T177 ,T178 ,T179 ,T180 ,T181 ,T182 ,T183 ,T184 ,T185 ,T186 ,T187 ,T188 ,T189 ,T190 ,T191 ,T192 ,T193 ,T194 ,T195 ,T196 ,T197 ,T198 ,T199 ,T200 ,T201;
wire 	 Z1 ,Z2 ,Z3 ,Z4 ,Z5 ,Z6 ,Z7 ,Z8 ,Z9 ,Z10 ,Z11 ,Z12 ,Z13 ,Z14 ,Z15 ,Z16 ,Z17 ,Z18 ,Z19 ,Z20 ,Z21 ,Z22 ,Z23 ,Z24 ,Z25 ,Z26 ,Z27 ,Z28 ,Z29 ,Z30 ,Z31 ,Z32 ,Z33 ,Z34 ,Z35 ,Z36 ,Z37 ,Z38 ,Z39 ,Z40 ,Z41 ,Z42 ,Z43 ,Z44 ,Z45 ,Z46 ,Z47 ,Z48 ,Z49 ,Z50 ,Z51 ,Z52 ,Z53 ,Z54 ,Z55 ,Z56 ,Z57 ,Z58 ,Z59 ,Z60 ,Z61 ,Z62 ,Z63 ,Z64 ,Z65 ,Z66 ,Z67 ,Z68 ,Z69 ,Z70 ,Z71 ,Z72 ,Z73 ,Z74 ,Z75 ,Z76 ,Z77 ,Z78 ,Z79 ,Z80 ,Z81 ,Z82 ,Z83 ,Z84 ,Z85 ,Z86 ,Z87 ,Z88 ,Z89 ,Z90 ,Z91 ,Z92 ,Z93 ,Z94 ,Z95 ,Z96 ,Z97 ,Z98 ,Z99 ,Z100 ,Z101 ,Z102 ,Z103 ,Z104 ,Z105 ,Z106 ,Z107 ,Z108 ,Z109 ,Z110 ,Z111 ,Z112 ,Z113 ,Z114 ,Z115 ,Z116 ,Z117 ,Z118 ,Z119 ,Z120 ,Z121 ,Z122 ,Z123 ,Z124 ,Z125 ,Z126 ,Z127 ,Z128 ,Z129 ,Z130 ,Z131 ,Z132 ,Z133 ,Z134 ,Z135 ,Z136 ,Z137 ,Z138 ,Z139 ,Z140 ,Z141 ,Z142 ,Z143 ,Z144 ,Z145 ,Z146 ,Z147 ,Z148 ,Z149 ,Z150 ,Z151 ,Z152 ,Z153 ,Z154 ,Z155 ,Z156 ,Z157 ,Z158 ,Z159 ,Z160 ,Z161 ,Z162 ,Z163 ,Z164 ,Z165 ,Z166 ,Z167 ,Z168 ,Z169 ,Z170 ,Z171 ,Z172 ,Z173 ,Z174 ,Z175 ,Z176 ,Z177 ,Z178 ,Z179 ,Z180 ,Z181 ,Z182 ,Z183 ,Z184 ,Z185 ,Z186 ,Z187 ,Z188 ,Z189 ,Z190 ,Z191 ,Z192 ,Z193 ,Z194 ,Z195 ,Z196 ,Z197 ,Z198 ,Z199 ,Z200;
medianCell_leftMst  m1(.X(X), .clk(clk), .reset(reset), .W(W), .isMedian(isLast1|isLast2), .R1_R(R1_2), .R_old_in(R_old), .T_R(T2), .R1(R1_1), .R2(R2_1), .R_median(median), .R_old_out(R_old), .Z(Z1), .T(T1), .isLast(isLast1));
medianFilterCell  m2(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd2), .isMedian(isLast3|isLast4), .R1_L(R1_1), .R1_R(R1_3), .R2_L(R2_1), .R_old_in(R_old), .Z_L(Z1), .T_L(T1), .T_R(T3), .R1(R1_2), .R2(R2_2), .R_median(median), .R_old_out(R_old), .Z(Z2), .T(T2), .isLast(isLast2));
medianFilterCell  m3(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd3), .isMedian(isLast5|isLast6), .R1_L(R1_2), .R1_R(R1_4), .R2_L(R2_2), .R_old_in(R_old), .Z_L(Z2), .T_L(T2), .T_R(T4), .R1(R1_3), .R2(R2_3), .R_median(median), .R_old_out(R_old), .Z(Z3), .T(T3), .isLast(isLast3));
medianFilterCell  m4(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd4), .isMedian(isLast7|isLast8), .R1_L(R1_3), .R1_R(R1_5), .R2_L(R2_3), .R_old_in(R_old), .Z_L(Z3), .T_L(T3), .T_R(T5), .R1(R1_4), .R2(R2_4), .R_median(median), .R_old_out(R_old), .Z(Z4), .T(T4), .isLast(isLast4));
medianFilterCell  m5(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd5), .isMedian(isLast9|isLast10), .R1_L(R1_4), .R1_R(R1_6), .R2_L(R2_4), .R_old_in(R_old), .Z_L(Z4), .T_L(T4), .T_R(T6), .R1(R1_5), .R2(R2_5), .R_median(median), .R_old_out(R_old), .Z(Z5), .T(T5), .isLast(isLast5));
medianFilterCell  m6(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd6), .isMedian(isLast11|isLast12), .R1_L(R1_5), .R1_R(R1_7), .R2_L(R2_5), .R_old_in(R_old), .Z_L(Z5), .T_L(T5), .T_R(T7), .R1(R1_6), .R2(R2_6), .R_median(median), .R_old_out(R_old), .Z(Z6), .T(T6), .isLast(isLast6));
medianFilterCell  m7(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd7), .isMedian(isLast13|isLast14), .R1_L(R1_6), .R1_R(R1_8), .R2_L(R2_6), .R_old_in(R_old), .Z_L(Z6), .T_L(T6), .T_R(T8), .R1(R1_7), .R2(R2_7), .R_median(median), .R_old_out(R_old), .Z(Z7), .T(T7), .isLast(isLast7));
medianFilterCell  m8(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd8), .isMedian(isLast15|isLast16), .R1_L(R1_7), .R1_R(R1_9), .R2_L(R2_7), .R_old_in(R_old), .Z_L(Z7), .T_L(T7), .T_R(T9), .R1(R1_8), .R2(R2_8), .R_median(median), .R_old_out(R_old), .Z(Z8), .T(T8), .isLast(isLast8));
medianFilterCell  m9(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd9), .isMedian(isLast17|isLast18), .R1_L(R1_8), .R1_R(R1_10), .R2_L(R2_8), .R_old_in(R_old), .Z_L(Z8), .T_L(T8), .T_R(T10), .R1(R1_9), .R2(R2_9), .R_median(median), .R_old_out(R_old), .Z(Z9), .T(T9), .isLast(isLast9));
medianFilterCell  m10(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd10), .isMedian(isLast19|isLast20), .R1_L(R1_9), .R1_R(R1_11), .R2_L(R2_9), .R_old_in(R_old), .Z_L(Z9), .T_L(T9), .T_R(T11), .R1(R1_10), .R2(R2_10), .R_median(median), .R_old_out(R_old), .Z(Z10), .T(T10), .isLast(isLast10));
medianFilterCell  m11(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd11), .isMedian(isLast21|isLast22), .R1_L(R1_10), .R1_R(R1_12), .R2_L(R2_10), .R_old_in(R_old), .Z_L(Z10), .T_L(T10), .T_R(T12), .R1(R1_11), .R2(R2_11), .R_median(median), .R_old_out(R_old), .Z(Z11), .T(T11), .isLast(isLast11));
medianFilterCell  m12(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd12), .isMedian(isLast23|isLast24), .R1_L(R1_11), .R1_R(R1_13), .R2_L(R2_11), .R_old_in(R_old), .Z_L(Z11), .T_L(T11), .T_R(T13), .R1(R1_12), .R2(R2_12), .R_median(median), .R_old_out(R_old), .Z(Z12), .T(T12), .isLast(isLast12));
medianFilterCell  m13(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd13), .isMedian(isLast25|isLast26), .R1_L(R1_12), .R1_R(R1_14), .R2_L(R2_12), .R_old_in(R_old), .Z_L(Z12), .T_L(T12), .T_R(T14), .R1(R1_13), .R2(R2_13), .R_median(median), .R_old_out(R_old), .Z(Z13), .T(T13), .isLast(isLast13));
medianFilterCell  m14(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd14), .isMedian(isLast27|isLast28), .R1_L(R1_13), .R1_R(R1_15), .R2_L(R2_13), .R_old_in(R_old), .Z_L(Z13), .T_L(T13), .T_R(T15), .R1(R1_14), .R2(R2_14), .R_median(median), .R_old_out(R_old), .Z(Z14), .T(T14), .isLast(isLast14));
medianFilterCell  m15(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd15), .isMedian(isLast29|isLast30), .R1_L(R1_14), .R1_R(R1_16), .R2_L(R2_14), .R_old_in(R_old), .Z_L(Z14), .T_L(T14), .T_R(T16), .R1(R1_15), .R2(R2_15), .R_median(median), .R_old_out(R_old), .Z(Z15), .T(T15), .isLast(isLast15));
medianFilterCell  m16(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd16), .isMedian(isLast31|isLast32), .R1_L(R1_15), .R1_R(R1_17), .R2_L(R2_15), .R_old_in(R_old), .Z_L(Z15), .T_L(T15), .T_R(T17), .R1(R1_16), .R2(R2_16), .R_median(median), .R_old_out(R_old), .Z(Z16), .T(T16), .isLast(isLast16));
medianFilterCell  m17(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd17), .isMedian(isLast33|isLast34), .R1_L(R1_16), .R1_R(R1_18), .R2_L(R2_16), .R_old_in(R_old), .Z_L(Z16), .T_L(T16), .T_R(T18), .R1(R1_17), .R2(R2_17), .R_median(median), .R_old_out(R_old), .Z(Z17), .T(T17), .isLast(isLast17));
medianFilterCell  m18(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd18), .isMedian(isLast35|isLast36), .R1_L(R1_17), .R1_R(R1_19), .R2_L(R2_17), .R_old_in(R_old), .Z_L(Z17), .T_L(T17), .T_R(T19), .R1(R1_18), .R2(R2_18), .R_median(median), .R_old_out(R_old), .Z(Z18), .T(T18), .isLast(isLast18));
medianFilterCell  m19(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd19), .isMedian(isLast37|isLast38), .R1_L(R1_18), .R1_R(R1_20), .R2_L(R2_18), .R_old_in(R_old), .Z_L(Z18), .T_L(T18), .T_R(T20), .R1(R1_19), .R2(R2_19), .R_median(median), .R_old_out(R_old), .Z(Z19), .T(T19), .isLast(isLast19));
medianFilterCell  m20(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd20), .isMedian(isLast39|isLast40), .R1_L(R1_19), .R1_R(R1_21), .R2_L(R2_19), .R_old_in(R_old), .Z_L(Z19), .T_L(T19), .T_R(T21), .R1(R1_20), .R2(R2_20), .R_median(median), .R_old_out(R_old), .Z(Z20), .T(T20), .isLast(isLast20));
medianFilterCell  m21(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd21), .isMedian(isLast41|isLast42), .R1_L(R1_20), .R1_R(R1_22), .R2_L(R2_20), .R_old_in(R_old), .Z_L(Z20), .T_L(T20), .T_R(T22), .R1(R1_21), .R2(R2_21), .R_median(median), .R_old_out(R_old), .Z(Z21), .T(T21), .isLast(isLast21));
medianFilterCell  m22(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd22), .isMedian(isLast43|isLast44), .R1_L(R1_21), .R1_R(R1_23), .R2_L(R2_21), .R_old_in(R_old), .Z_L(Z21), .T_L(T21), .T_R(T23), .R1(R1_22), .R2(R2_22), .R_median(median), .R_old_out(R_old), .Z(Z22), .T(T22), .isLast(isLast22));
medianFilterCell  m23(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd23), .isMedian(isLast45|isLast46), .R1_L(R1_22), .R1_R(R1_24), .R2_L(R2_22), .R_old_in(R_old), .Z_L(Z22), .T_L(T22), .T_R(T24), .R1(R1_23), .R2(R2_23), .R_median(median), .R_old_out(R_old), .Z(Z23), .T(T23), .isLast(isLast23));
medianFilterCell  m24(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd24), .isMedian(isLast47|isLast48), .R1_L(R1_23), .R1_R(R1_25), .R2_L(R2_23), .R_old_in(R_old), .Z_L(Z23), .T_L(T23), .T_R(T25), .R1(R1_24), .R2(R2_24), .R_median(median), .R_old_out(R_old), .Z(Z24), .T(T24), .isLast(isLast24));
medianFilterCell  m25(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd25), .isMedian(isLast49|isLast50), .R1_L(R1_24), .R1_R(R1_26), .R2_L(R2_24), .R_old_in(R_old), .Z_L(Z24), .T_L(T24), .T_R(T26), .R1(R1_25), .R2(R2_25), .R_median(median), .R_old_out(R_old), .Z(Z25), .T(T25), .isLast(isLast25));
medianFilterCell  m26(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd26), .isMedian(isLast51|isLast52), .R1_L(R1_25), .R1_R(R1_27), .R2_L(R2_25), .R_old_in(R_old), .Z_L(Z25), .T_L(T25), .T_R(T27), .R1(R1_26), .R2(R2_26), .R_median(median), .R_old_out(R_old), .Z(Z26), .T(T26), .isLast(isLast26));
medianFilterCell  m27(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd27), .isMedian(isLast53|isLast54), .R1_L(R1_26), .R1_R(R1_28), .R2_L(R2_26), .R_old_in(R_old), .Z_L(Z26), .T_L(T26), .T_R(T28), .R1(R1_27), .R2(R2_27), .R_median(median), .R_old_out(R_old), .Z(Z27), .T(T27), .isLast(isLast27));
medianFilterCell  m28(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd28), .isMedian(isLast55|isLast56), .R1_L(R1_27), .R1_R(R1_29), .R2_L(R2_27), .R_old_in(R_old), .Z_L(Z27), .T_L(T27), .T_R(T29), .R1(R1_28), .R2(R2_28), .R_median(median), .R_old_out(R_old), .Z(Z28), .T(T28), .isLast(isLast28));
medianFilterCell  m29(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd29), .isMedian(isLast57|isLast58), .R1_L(R1_28), .R1_R(R1_30), .R2_L(R2_28), .R_old_in(R_old), .Z_L(Z28), .T_L(T28), .T_R(T30), .R1(R1_29), .R2(R2_29), .R_median(median), .R_old_out(R_old), .Z(Z29), .T(T29), .isLast(isLast29));
medianFilterCell  m30(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd30), .isMedian(isLast59|isLast60), .R1_L(R1_29), .R1_R(R1_31), .R2_L(R2_29), .R_old_in(R_old), .Z_L(Z29), .T_L(T29), .T_R(T31), .R1(R1_30), .R2(R2_30), .R_median(median), .R_old_out(R_old), .Z(Z30), .T(T30), .isLast(isLast30));
medianFilterCell  m31(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd31), .isMedian(isLast61|isLast62), .R1_L(R1_30), .R1_R(R1_32), .R2_L(R2_30), .R_old_in(R_old), .Z_L(Z30), .T_L(T30), .T_R(T32), .R1(R1_31), .R2(R2_31), .R_median(median), .R_old_out(R_old), .Z(Z31), .T(T31), .isLast(isLast31));
medianFilterCell  m32(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd32), .isMedian(isLast63|isLast64), .R1_L(R1_31), .R1_R(R1_33), .R2_L(R2_31), .R_old_in(R_old), .Z_L(Z31), .T_L(T31), .T_R(T33), .R1(R1_32), .R2(R2_32), .R_median(median), .R_old_out(R_old), .Z(Z32), .T(T32), .isLast(isLast32));
medianFilterCell  m33(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd33), .isMedian(isLast65|isLast66), .R1_L(R1_32), .R1_R(R1_34), .R2_L(R2_32), .R_old_in(R_old), .Z_L(Z32), .T_L(T32), .T_R(T34), .R1(R1_33), .R2(R2_33), .R_median(median), .R_old_out(R_old), .Z(Z33), .T(T33), .isLast(isLast33));
medianFilterCell  m34(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd34), .isMedian(isLast67|isLast68), .R1_L(R1_33), .R1_R(R1_35), .R2_L(R2_33), .R_old_in(R_old), .Z_L(Z33), .T_L(T33), .T_R(T35), .R1(R1_34), .R2(R2_34), .R_median(median), .R_old_out(R_old), .Z(Z34), .T(T34), .isLast(isLast34));
medianFilterCell  m35(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd35), .isMedian(isLast69|isLast70), .R1_L(R1_34), .R1_R(R1_36), .R2_L(R2_34), .R_old_in(R_old), .Z_L(Z34), .T_L(T34), .T_R(T36), .R1(R1_35), .R2(R2_35), .R_median(median), .R_old_out(R_old), .Z(Z35), .T(T35), .isLast(isLast35));
medianFilterCell  m36(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd36), .isMedian(isLast71|isLast72), .R1_L(R1_35), .R1_R(R1_37), .R2_L(R2_35), .R_old_in(R_old), .Z_L(Z35), .T_L(T35), .T_R(T37), .R1(R1_36), .R2(R2_36), .R_median(median), .R_old_out(R_old), .Z(Z36), .T(T36), .isLast(isLast36));
medianFilterCell  m37(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd37), .isMedian(isLast73|isLast74), .R1_L(R1_36), .R1_R(R1_38), .R2_L(R2_36), .R_old_in(R_old), .Z_L(Z36), .T_L(T36), .T_R(T38), .R1(R1_37), .R2(R2_37), .R_median(median), .R_old_out(R_old), .Z(Z37), .T(T37), .isLast(isLast37));
medianFilterCell  m38(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd38), .isMedian(isLast75|isLast76), .R1_L(R1_37), .R1_R(R1_39), .R2_L(R2_37), .R_old_in(R_old), .Z_L(Z37), .T_L(T37), .T_R(T39), .R1(R1_38), .R2(R2_38), .R_median(median), .R_old_out(R_old), .Z(Z38), .T(T38), .isLast(isLast38));
medianFilterCell  m39(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd39), .isMedian(isLast77|isLast78), .R1_L(R1_38), .R1_R(R1_40), .R2_L(R2_38), .R_old_in(R_old), .Z_L(Z38), .T_L(T38), .T_R(T40), .R1(R1_39), .R2(R2_39), .R_median(median), .R_old_out(R_old), .Z(Z39), .T(T39), .isLast(isLast39));
medianFilterCell  m40(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd40), .isMedian(isLast79|isLast80), .R1_L(R1_39), .R1_R(R1_41), .R2_L(R2_39), .R_old_in(R_old), .Z_L(Z39), .T_L(T39), .T_R(T41), .R1(R1_40), .R2(R2_40), .R_median(median), .R_old_out(R_old), .Z(Z40), .T(T40), .isLast(isLast40));
medianFilterCell  m41(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd41), .isMedian(isLast81|isLast82), .R1_L(R1_40), .R1_R(R1_42), .R2_L(R2_40), .R_old_in(R_old), .Z_L(Z40), .T_L(T40), .T_R(T42), .R1(R1_41), .R2(R2_41), .R_median(median), .R_old_out(R_old), .Z(Z41), .T(T41), .isLast(isLast41));
medianFilterCell  m42(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd42), .isMedian(isLast83|isLast84), .R1_L(R1_41), .R1_R(R1_43), .R2_L(R2_41), .R_old_in(R_old), .Z_L(Z41), .T_L(T41), .T_R(T43), .R1(R1_42), .R2(R2_42), .R_median(median), .R_old_out(R_old), .Z(Z42), .T(T42), .isLast(isLast42));
medianFilterCell  m43(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd43), .isMedian(isLast85|isLast86), .R1_L(R1_42), .R1_R(R1_44), .R2_L(R2_42), .R_old_in(R_old), .Z_L(Z42), .T_L(T42), .T_R(T44), .R1(R1_43), .R2(R2_43), .R_median(median), .R_old_out(R_old), .Z(Z43), .T(T43), .isLast(isLast43));
medianFilterCell  m44(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd44), .isMedian(isLast87|isLast88), .R1_L(R1_43), .R1_R(R1_45), .R2_L(R2_43), .R_old_in(R_old), .Z_L(Z43), .T_L(T43), .T_R(T45), .R1(R1_44), .R2(R2_44), .R_median(median), .R_old_out(R_old), .Z(Z44), .T(T44), .isLast(isLast44));
medianFilterCell  m45(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd45), .isMedian(isLast89|isLast90), .R1_L(R1_44), .R1_R(R1_46), .R2_L(R2_44), .R_old_in(R_old), .Z_L(Z44), .T_L(T44), .T_R(T46), .R1(R1_45), .R2(R2_45), .R_median(median), .R_old_out(R_old), .Z(Z45), .T(T45), .isLast(isLast45));
medianFilterCell  m46(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd46), .isMedian(isLast91|isLast92), .R1_L(R1_45), .R1_R(R1_47), .R2_L(R2_45), .R_old_in(R_old), .Z_L(Z45), .T_L(T45), .T_R(T47), .R1(R1_46), .R2(R2_46), .R_median(median), .R_old_out(R_old), .Z(Z46), .T(T46), .isLast(isLast46));
medianFilterCell  m47(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd47), .isMedian(isLast93|isLast94), .R1_L(R1_46), .R1_R(R1_48), .R2_L(R2_46), .R_old_in(R_old), .Z_L(Z46), .T_L(T46), .T_R(T48), .R1(R1_47), .R2(R2_47), .R_median(median), .R_old_out(R_old), .Z(Z47), .T(T47), .isLast(isLast47));
medianFilterCell  m48(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd48), .isMedian(isLast95|isLast96), .R1_L(R1_47), .R1_R(R1_49), .R2_L(R2_47), .R_old_in(R_old), .Z_L(Z47), .T_L(T47), .T_R(T49), .R1(R1_48), .R2(R2_48), .R_median(median), .R_old_out(R_old), .Z(Z48), .T(T48), .isLast(isLast48));
medianFilterCell  m49(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd49), .isMedian(isLast97|isLast98), .R1_L(R1_48), .R1_R(R1_50), .R2_L(R2_48), .R_old_in(R_old), .Z_L(Z48), .T_L(T48), .T_R(T50), .R1(R1_49), .R2(R2_49), .R_median(median), .R_old_out(R_old), .Z(Z49), .T(T49), .isLast(isLast49));
medianFilterCell  m50(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd50), .isMedian(isLast99|isLast100), .R1_L(R1_49), .R1_R(R1_51), .R2_L(R2_49), .R_old_in(R_old), .Z_L(Z49), .T_L(T49), .T_R(T51), .R1(R1_50), .R2(R2_50), .R_median(median), .R_old_out(R_old), .Z(Z50), .T(T50), .isLast(isLast50));
medianFilterCell  m51(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd51), .isMedian(isLast101|isLast102), .R1_L(R1_50), .R1_R(R1_52), .R2_L(R2_50), .R_old_in(R_old), .Z_L(Z50), .T_L(T50), .T_R(T52), .R1(R1_51), .R2(R2_51), .R_median(median), .R_old_out(R_old), .Z(Z51), .T(T51), .isLast(isLast51));
medianFilterCell  m52(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd52), .isMedian(isLast103|isLast104), .R1_L(R1_51), .R1_R(R1_53), .R2_L(R2_51), .R_old_in(R_old), .Z_L(Z51), .T_L(T51), .T_R(T53), .R1(R1_52), .R2(R2_52), .R_median(median), .R_old_out(R_old), .Z(Z52), .T(T52), .isLast(isLast52));
medianFilterCell  m53(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd53), .isMedian(isLast105|isLast106), .R1_L(R1_52), .R1_R(R1_54), .R2_L(R2_52), .R_old_in(R_old), .Z_L(Z52), .T_L(T52), .T_R(T54), .R1(R1_53), .R2(R2_53), .R_median(median), .R_old_out(R_old), .Z(Z53), .T(T53), .isLast(isLast53));
medianFilterCell  m54(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd54), .isMedian(isLast107|isLast108), .R1_L(R1_53), .R1_R(R1_55), .R2_L(R2_53), .R_old_in(R_old), .Z_L(Z53), .T_L(T53), .T_R(T55), .R1(R1_54), .R2(R2_54), .R_median(median), .R_old_out(R_old), .Z(Z54), .T(T54), .isLast(isLast54));
medianFilterCell  m55(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd55), .isMedian(isLast109|isLast110), .R1_L(R1_54), .R1_R(R1_56), .R2_L(R2_54), .R_old_in(R_old), .Z_L(Z54), .T_L(T54), .T_R(T56), .R1(R1_55), .R2(R2_55), .R_median(median), .R_old_out(R_old), .Z(Z55), .T(T55), .isLast(isLast55));
medianFilterCell  m56(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd56), .isMedian(isLast111|isLast112), .R1_L(R1_55), .R1_R(R1_57), .R2_L(R2_55), .R_old_in(R_old), .Z_L(Z55), .T_L(T55), .T_R(T57), .R1(R1_56), .R2(R2_56), .R_median(median), .R_old_out(R_old), .Z(Z56), .T(T56), .isLast(isLast56));
medianFilterCell  m57(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd57), .isMedian(isLast113|isLast114), .R1_L(R1_56), .R1_R(R1_58), .R2_L(R2_56), .R_old_in(R_old), .Z_L(Z56), .T_L(T56), .T_R(T58), .R1(R1_57), .R2(R2_57), .R_median(median), .R_old_out(R_old), .Z(Z57), .T(T57), .isLast(isLast57));
medianFilterCell  m58(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd58), .isMedian(isLast115|isLast116), .R1_L(R1_57), .R1_R(R1_59), .R2_L(R2_57), .R_old_in(R_old), .Z_L(Z57), .T_L(T57), .T_R(T59), .R1(R1_58), .R2(R2_58), .R_median(median), .R_old_out(R_old), .Z(Z58), .T(T58), .isLast(isLast58));
medianFilterCell  m59(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd59), .isMedian(isLast117|isLast118), .R1_L(R1_58), .R1_R(R1_60), .R2_L(R2_58), .R_old_in(R_old), .Z_L(Z58), .T_L(T58), .T_R(T60), .R1(R1_59), .R2(R2_59), .R_median(median), .R_old_out(R_old), .Z(Z59), .T(T59), .isLast(isLast59));
medianFilterCell  m60(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd60), .isMedian(isLast119|isLast120), .R1_L(R1_59), .R1_R(R1_61), .R2_L(R2_59), .R_old_in(R_old), .Z_L(Z59), .T_L(T59), .T_R(T61), .R1(R1_60), .R2(R2_60), .R_median(median), .R_old_out(R_old), .Z(Z60), .T(T60), .isLast(isLast60));
medianFilterCell  m61(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd61), .isMedian(isLast121|isLast122), .R1_L(R1_60), .R1_R(R1_62), .R2_L(R2_60), .R_old_in(R_old), .Z_L(Z60), .T_L(T60), .T_R(T62), .R1(R1_61), .R2(R2_61), .R_median(median), .R_old_out(R_old), .Z(Z61), .T(T61), .isLast(isLast61));
medianFilterCell  m62(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd62), .isMedian(isLast123|isLast124), .R1_L(R1_61), .R1_R(R1_63), .R2_L(R2_61), .R_old_in(R_old), .Z_L(Z61), .T_L(T61), .T_R(T63), .R1(R1_62), .R2(R2_62), .R_median(median), .R_old_out(R_old), .Z(Z62), .T(T62), .isLast(isLast62));
medianFilterCell  m63(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd63), .isMedian(isLast125|isLast126), .R1_L(R1_62), .R1_R(R1_64), .R2_L(R2_62), .R_old_in(R_old), .Z_L(Z62), .T_L(T62), .T_R(T64), .R1(R1_63), .R2(R2_63), .R_median(median), .R_old_out(R_old), .Z(Z63), .T(T63), .isLast(isLast63));
medianFilterCell  m64(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd64), .isMedian(isLast127|isLast128), .R1_L(R1_63), .R1_R(R1_65), .R2_L(R2_63), .R_old_in(R_old), .Z_L(Z63), .T_L(T63), .T_R(T65), .R1(R1_64), .R2(R2_64), .R_median(median), .R_old_out(R_old), .Z(Z64), .T(T64), .isLast(isLast64));
medianFilterCell  m65(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd65), .isMedian(isLast129|isLast130), .R1_L(R1_64), .R1_R(R1_66), .R2_L(R2_64), .R_old_in(R_old), .Z_L(Z64), .T_L(T64), .T_R(T66), .R1(R1_65), .R2(R2_65), .R_median(median), .R_old_out(R_old), .Z(Z65), .T(T65), .isLast(isLast65));
medianFilterCell  m66(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd66), .isMedian(isLast131|isLast132), .R1_L(R1_65), .R1_R(R1_67), .R2_L(R2_65), .R_old_in(R_old), .Z_L(Z65), .T_L(T65), .T_R(T67), .R1(R1_66), .R2(R2_66), .R_median(median), .R_old_out(R_old), .Z(Z66), .T(T66), .isLast(isLast66));
medianFilterCell  m67(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd67), .isMedian(isLast133|isLast134), .R1_L(R1_66), .R1_R(R1_68), .R2_L(R2_66), .R_old_in(R_old), .Z_L(Z66), .T_L(T66), .T_R(T68), .R1(R1_67), .R2(R2_67), .R_median(median), .R_old_out(R_old), .Z(Z67), .T(T67), .isLast(isLast67));
medianFilterCell  m68(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd68), .isMedian(isLast135|isLast136), .R1_L(R1_67), .R1_R(R1_69), .R2_L(R2_67), .R_old_in(R_old), .Z_L(Z67), .T_L(T67), .T_R(T69), .R1(R1_68), .R2(R2_68), .R_median(median), .R_old_out(R_old), .Z(Z68), .T(T68), .isLast(isLast68));
medianFilterCell  m69(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd69), .isMedian(isLast137|isLast138), .R1_L(R1_68), .R1_R(R1_70), .R2_L(R2_68), .R_old_in(R_old), .Z_L(Z68), .T_L(T68), .T_R(T70), .R1(R1_69), .R2(R2_69), .R_median(median), .R_old_out(R_old), .Z(Z69), .T(T69), .isLast(isLast69));
medianFilterCell  m70(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd70), .isMedian(isLast139|isLast140), .R1_L(R1_69), .R1_R(R1_71), .R2_L(R2_69), .R_old_in(R_old), .Z_L(Z69), .T_L(T69), .T_R(T71), .R1(R1_70), .R2(R2_70), .R_median(median), .R_old_out(R_old), .Z(Z70), .T(T70), .isLast(isLast70));
medianFilterCell  m71(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd71), .isMedian(isLast141|isLast142), .R1_L(R1_70), .R1_R(R1_72), .R2_L(R2_70), .R_old_in(R_old), .Z_L(Z70), .T_L(T70), .T_R(T72), .R1(R1_71), .R2(R2_71), .R_median(median), .R_old_out(R_old), .Z(Z71), .T(T71), .isLast(isLast71));
medianFilterCell  m72(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd72), .isMedian(isLast143|isLast144), .R1_L(R1_71), .R1_R(R1_73), .R2_L(R2_71), .R_old_in(R_old), .Z_L(Z71), .T_L(T71), .T_R(T73), .R1(R1_72), .R2(R2_72), .R_median(median), .R_old_out(R_old), .Z(Z72), .T(T72), .isLast(isLast72));
medianFilterCell  m73(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd73), .isMedian(isLast145|isLast146), .R1_L(R1_72), .R1_R(R1_74), .R2_L(R2_72), .R_old_in(R_old), .Z_L(Z72), .T_L(T72), .T_R(T74), .R1(R1_73), .R2(R2_73), .R_median(median), .R_old_out(R_old), .Z(Z73), .T(T73), .isLast(isLast73));
medianFilterCell  m74(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd74), .isMedian(isLast147|isLast148), .R1_L(R1_73), .R1_R(R1_75), .R2_L(R2_73), .R_old_in(R_old), .Z_L(Z73), .T_L(T73), .T_R(T75), .R1(R1_74), .R2(R2_74), .R_median(median), .R_old_out(R_old), .Z(Z74), .T(T74), .isLast(isLast74));
medianFilterCell  m75(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd75), .isMedian(isLast149|isLast150), .R1_L(R1_74), .R1_R(R1_76), .R2_L(R2_74), .R_old_in(R_old), .Z_L(Z74), .T_L(T74), .T_R(T76), .R1(R1_75), .R2(R2_75), .R_median(median), .R_old_out(R_old), .Z(Z75), .T(T75), .isLast(isLast75));
medianFilterCell  m76(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd76), .isMedian(isLast151|isLast152), .R1_L(R1_75), .R1_R(R1_77), .R2_L(R2_75), .R_old_in(R_old), .Z_L(Z75), .T_L(T75), .T_R(T77), .R1(R1_76), .R2(R2_76), .R_median(median), .R_old_out(R_old), .Z(Z76), .T(T76), .isLast(isLast76));
medianFilterCell  m77(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd77), .isMedian(isLast153|isLast154), .R1_L(R1_76), .R1_R(R1_78), .R2_L(R2_76), .R_old_in(R_old), .Z_L(Z76), .T_L(T76), .T_R(T78), .R1(R1_77), .R2(R2_77), .R_median(median), .R_old_out(R_old), .Z(Z77), .T(T77), .isLast(isLast77));
medianFilterCell  m78(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd78), .isMedian(isLast155|isLast156), .R1_L(R1_77), .R1_R(R1_79), .R2_L(R2_77), .R_old_in(R_old), .Z_L(Z77), .T_L(T77), .T_R(T79), .R1(R1_78), .R2(R2_78), .R_median(median), .R_old_out(R_old), .Z(Z78), .T(T78), .isLast(isLast78));
medianFilterCell  m79(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd79), .isMedian(isLast157|isLast158), .R1_L(R1_78), .R1_R(R1_80), .R2_L(R2_78), .R_old_in(R_old), .Z_L(Z78), .T_L(T78), .T_R(T80), .R1(R1_79), .R2(R2_79), .R_median(median), .R_old_out(R_old), .Z(Z79), .T(T79), .isLast(isLast79));
medianFilterCell  m80(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd80), .isMedian(isLast159|isLast160), .R1_L(R1_79), .R1_R(R1_81), .R2_L(R2_79), .R_old_in(R_old), .Z_L(Z79), .T_L(T79), .T_R(T81), .R1(R1_80), .R2(R2_80), .R_median(median), .R_old_out(R_old), .Z(Z80), .T(T80), .isLast(isLast80));
medianFilterCell  m81(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd81), .isMedian(isLast161|isLast162), .R1_L(R1_80), .R1_R(R1_82), .R2_L(R2_80), .R_old_in(R_old), .Z_L(Z80), .T_L(T80), .T_R(T82), .R1(R1_81), .R2(R2_81), .R_median(median), .R_old_out(R_old), .Z(Z81), .T(T81), .isLast(isLast81));
medianFilterCell  m82(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd82), .isMedian(isLast163|isLast164), .R1_L(R1_81), .R1_R(R1_83), .R2_L(R2_81), .R_old_in(R_old), .Z_L(Z81), .T_L(T81), .T_R(T83), .R1(R1_82), .R2(R2_82), .R_median(median), .R_old_out(R_old), .Z(Z82), .T(T82), .isLast(isLast82));
medianFilterCell  m83(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd83), .isMedian(isLast165|isLast166), .R1_L(R1_82), .R1_R(R1_84), .R2_L(R2_82), .R_old_in(R_old), .Z_L(Z82), .T_L(T82), .T_R(T84), .R1(R1_83), .R2(R2_83), .R_median(median), .R_old_out(R_old), .Z(Z83), .T(T83), .isLast(isLast83));
medianFilterCell  m84(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd84), .isMedian(isLast167|isLast168), .R1_L(R1_83), .R1_R(R1_85), .R2_L(R2_83), .R_old_in(R_old), .Z_L(Z83), .T_L(T83), .T_R(T85), .R1(R1_84), .R2(R2_84), .R_median(median), .R_old_out(R_old), .Z(Z84), .T(T84), .isLast(isLast84));
medianFilterCell  m85(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd85), .isMedian(isLast169|isLast170), .R1_L(R1_84), .R1_R(R1_86), .R2_L(R2_84), .R_old_in(R_old), .Z_L(Z84), .T_L(T84), .T_R(T86), .R1(R1_85), .R2(R2_85), .R_median(median), .R_old_out(R_old), .Z(Z85), .T(T85), .isLast(isLast85));
medianFilterCell  m86(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd86), .isMedian(isLast171|isLast172), .R1_L(R1_85), .R1_R(R1_87), .R2_L(R2_85), .R_old_in(R_old), .Z_L(Z85), .T_L(T85), .T_R(T87), .R1(R1_86), .R2(R2_86), .R_median(median), .R_old_out(R_old), .Z(Z86), .T(T86), .isLast(isLast86));
medianFilterCell  m87(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd87), .isMedian(isLast173|isLast174), .R1_L(R1_86), .R1_R(R1_88), .R2_L(R2_86), .R_old_in(R_old), .Z_L(Z86), .T_L(T86), .T_R(T88), .R1(R1_87), .R2(R2_87), .R_median(median), .R_old_out(R_old), .Z(Z87), .T(T87), .isLast(isLast87));
medianFilterCell  m88(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd88), .isMedian(isLast175|isLast176), .R1_L(R1_87), .R1_R(R1_89), .R2_L(R2_87), .R_old_in(R_old), .Z_L(Z87), .T_L(T87), .T_R(T89), .R1(R1_88), .R2(R2_88), .R_median(median), .R_old_out(R_old), .Z(Z88), .T(T88), .isLast(isLast88));
medianFilterCell  m89(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd89), .isMedian(isLast177|isLast178), .R1_L(R1_88), .R1_R(R1_90), .R2_L(R2_88), .R_old_in(R_old), .Z_L(Z88), .T_L(T88), .T_R(T90), .R1(R1_89), .R2(R2_89), .R_median(median), .R_old_out(R_old), .Z(Z89), .T(T89), .isLast(isLast89));
medianFilterCell  m90(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd90), .isMedian(isLast179|isLast180), .R1_L(R1_89), .R1_R(R1_91), .R2_L(R2_89), .R_old_in(R_old), .Z_L(Z89), .T_L(T89), .T_R(T91), .R1(R1_90), .R2(R2_90), .R_median(median), .R_old_out(R_old), .Z(Z90), .T(T90), .isLast(isLast90));
medianFilterCell  m91(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd91), .isMedian(isLast181|isLast182), .R1_L(R1_90), .R1_R(R1_92), .R2_L(R2_90), .R_old_in(R_old), .Z_L(Z90), .T_L(T90), .T_R(T92), .R1(R1_91), .R2(R2_91), .R_median(median), .R_old_out(R_old), .Z(Z91), .T(T91), .isLast(isLast91));
medianFilterCell  m92(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd92), .isMedian(isLast183|isLast184), .R1_L(R1_91), .R1_R(R1_93), .R2_L(R2_91), .R_old_in(R_old), .Z_L(Z91), .T_L(T91), .T_R(T93), .R1(R1_92), .R2(R2_92), .R_median(median), .R_old_out(R_old), .Z(Z92), .T(T92), .isLast(isLast92));
medianFilterCell  m93(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd93), .isMedian(isLast185|isLast186), .R1_L(R1_92), .R1_R(R1_94), .R2_L(R2_92), .R_old_in(R_old), .Z_L(Z92), .T_L(T92), .T_R(T94), .R1(R1_93), .R2(R2_93), .R_median(median), .R_old_out(R_old), .Z(Z93), .T(T93), .isLast(isLast93));
medianFilterCell  m94(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd94), .isMedian(isLast187|isLast188), .R1_L(R1_93), .R1_R(R1_95), .R2_L(R2_93), .R_old_in(R_old), .Z_L(Z93), .T_L(T93), .T_R(T95), .R1(R1_94), .R2(R2_94), .R_median(median), .R_old_out(R_old), .Z(Z94), .T(T94), .isLast(isLast94));
medianFilterCell  m95(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd95), .isMedian(isLast189|isLast190), .R1_L(R1_94), .R1_R(R1_96), .R2_L(R2_94), .R_old_in(R_old), .Z_L(Z94), .T_L(T94), .T_R(T96), .R1(R1_95), .R2(R2_95), .R_median(median), .R_old_out(R_old), .Z(Z95), .T(T95), .isLast(isLast95));
medianFilterCell  m96(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd96), .isMedian(isLast191|isLast192), .R1_L(R1_95), .R1_R(R1_97), .R2_L(R2_95), .R_old_in(R_old), .Z_L(Z95), .T_L(T95), .T_R(T97), .R1(R1_96), .R2(R2_96), .R_median(median), .R_old_out(R_old), .Z(Z96), .T(T96), .isLast(isLast96));
medianFilterCell  m97(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd97), .isMedian(isLast193|isLast194), .R1_L(R1_96), .R1_R(R1_98), .R2_L(R2_96), .R_old_in(R_old), .Z_L(Z96), .T_L(T96), .T_R(T98), .R1(R1_97), .R2(R2_97), .R_median(median), .R_old_out(R_old), .Z(Z97), .T(T97), .isLast(isLast97));
medianFilterCell  m98(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd98), .isMedian(isLast195|isLast196), .R1_L(R1_97), .R1_R(R1_99), .R2_L(R2_97), .R_old_in(R_old), .Z_L(Z97), .T_L(T97), .T_R(T99), .R1(R1_98), .R2(R2_98), .R_median(median), .R_old_out(R_old), .Z(Z98), .T(T98), .isLast(isLast98));
medianFilterCell  m99(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd99), .isMedian(isLast197|isLast198), .R1_L(R1_98), .R1_R(R1_100), .R2_L(R2_98), .R_old_in(R_old), .Z_L(Z98), .T_L(T98), .T_R(T100), .R1(R1_99), .R2(R2_99), .R_median(median), .R_old_out(R_old), .Z(Z99), .T(T99), .isLast(isLast99));
medianFilterCell  m100(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd100), .isMedian(isLast199|isLast200), .R1_L(R1_99), .R1_R(R1_101), .R2_L(R2_99), .R_old_in(R_old), .Z_L(Z99), .T_L(T99), .T_R(T101), .R1(R1_100), .R2(R2_100), .R_median(median), .R_old_out(R_old), .Z(Z100), .T(T100), .isLast(isLast100));
medianFilterCell  m101(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd101), .isMedian(isLast201), .R1_L(R1_100), .R1_R(R1_102), .R2_L(R2_100), .R_old_in(R_old), .Z_L(Z100), .T_L(T100), .T_R(T102), .R1(R1_101), .R2(R2_101), .R_median(median), .R_old_out(R_old), .Z(Z101), .T(T101), .isLast(isLast101));
medianFilterCell  m102(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd102), .isMedian(1'b0), .R1_L(R1_101), .R1_R(R1_103), .R2_L(R2_101), .R_old_in(R_old), .Z_L(Z101), .T_L(T101), .T_R(T103), .R1(R1_102), .R2(R2_102), .R_median(median), .R_old_out(R_old), .Z(Z102), .T(T102), .isLast(isLast102));
medianFilterCell  m103(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd103), .isMedian(1'b0), .R1_L(R1_102), .R1_R(R1_104), .R2_L(R2_102), .R_old_in(R_old), .Z_L(Z102), .T_L(T102), .T_R(T104), .R1(R1_103), .R2(R2_103), .R_median(median), .R_old_out(R_old), .Z(Z103), .T(T103), .isLast(isLast103));
medianFilterCell  m104(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd104), .isMedian(1'b0), .R1_L(R1_103), .R1_R(R1_105), .R2_L(R2_103), .R_old_in(R_old), .Z_L(Z103), .T_L(T103), .T_R(T105), .R1(R1_104), .R2(R2_104), .R_median(median), .R_old_out(R_old), .Z(Z104), .T(T104), .isLast(isLast104));
medianFilterCell  m105(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd105), .isMedian(1'b0), .R1_L(R1_104), .R1_R(R1_106), .R2_L(R2_104), .R_old_in(R_old), .Z_L(Z104), .T_L(T104), .T_R(T106), .R1(R1_105), .R2(R2_105), .R_median(median), .R_old_out(R_old), .Z(Z105), .T(T105), .isLast(isLast105));
medianFilterCell  m106(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd106), .isMedian(1'b0), .R1_L(R1_105), .R1_R(R1_107), .R2_L(R2_105), .R_old_in(R_old), .Z_L(Z105), .T_L(T105), .T_R(T107), .R1(R1_106), .R2(R2_106), .R_median(median), .R_old_out(R_old), .Z(Z106), .T(T106), .isLast(isLast106));
medianFilterCell  m107(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd107), .isMedian(1'b0), .R1_L(R1_106), .R1_R(R1_108), .R2_L(R2_106), .R_old_in(R_old), .Z_L(Z106), .T_L(T106), .T_R(T108), .R1(R1_107), .R2(R2_107), .R_median(median), .R_old_out(R_old), .Z(Z107), .T(T107), .isLast(isLast107));
medianFilterCell  m108(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd108), .isMedian(1'b0), .R1_L(R1_107), .R1_R(R1_109), .R2_L(R2_107), .R_old_in(R_old), .Z_L(Z107), .T_L(T107), .T_R(T109), .R1(R1_108), .R2(R2_108), .R_median(median), .R_old_out(R_old), .Z(Z108), .T(T108), .isLast(isLast108));
medianFilterCell  m109(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd109), .isMedian(1'b0), .R1_L(R1_108), .R1_R(R1_110), .R2_L(R2_108), .R_old_in(R_old), .Z_L(Z108), .T_L(T108), .T_R(T110), .R1(R1_109), .R2(R2_109), .R_median(median), .R_old_out(R_old), .Z(Z109), .T(T109), .isLast(isLast109));
medianFilterCell  m110(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd110), .isMedian(1'b0), .R1_L(R1_109), .R1_R(R1_111), .R2_L(R2_109), .R_old_in(R_old), .Z_L(Z109), .T_L(T109), .T_R(T111), .R1(R1_110), .R2(R2_110), .R_median(median), .R_old_out(R_old), .Z(Z110), .T(T110), .isLast(isLast110));
medianFilterCell  m111(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd111), .isMedian(1'b0), .R1_L(R1_110), .R1_R(R1_112), .R2_L(R2_110), .R_old_in(R_old), .Z_L(Z110), .T_L(T110), .T_R(T112), .R1(R1_111), .R2(R2_111), .R_median(median), .R_old_out(R_old), .Z(Z111), .T(T111), .isLast(isLast111));
medianFilterCell  m112(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd112), .isMedian(1'b0), .R1_L(R1_111), .R1_R(R1_113), .R2_L(R2_111), .R_old_in(R_old), .Z_L(Z111), .T_L(T111), .T_R(T113), .R1(R1_112), .R2(R2_112), .R_median(median), .R_old_out(R_old), .Z(Z112), .T(T112), .isLast(isLast112));
medianFilterCell  m113(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd113), .isMedian(1'b0), .R1_L(R1_112), .R1_R(R1_114), .R2_L(R2_112), .R_old_in(R_old), .Z_L(Z112), .T_L(T112), .T_R(T114), .R1(R1_113), .R2(R2_113), .R_median(median), .R_old_out(R_old), .Z(Z113), .T(T113), .isLast(isLast113));
medianFilterCell  m114(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd114), .isMedian(1'b0), .R1_L(R1_113), .R1_R(R1_115), .R2_L(R2_113), .R_old_in(R_old), .Z_L(Z113), .T_L(T113), .T_R(T115), .R1(R1_114), .R2(R2_114), .R_median(median), .R_old_out(R_old), .Z(Z114), .T(T114), .isLast(isLast114));
medianFilterCell  m115(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd115), .isMedian(1'b0), .R1_L(R1_114), .R1_R(R1_116), .R2_L(R2_114), .R_old_in(R_old), .Z_L(Z114), .T_L(T114), .T_R(T116), .R1(R1_115), .R2(R2_115), .R_median(median), .R_old_out(R_old), .Z(Z115), .T(T115), .isLast(isLast115));
medianFilterCell  m116(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd116), .isMedian(1'b0), .R1_L(R1_115), .R1_R(R1_117), .R2_L(R2_115), .R_old_in(R_old), .Z_L(Z115), .T_L(T115), .T_R(T117), .R1(R1_116), .R2(R2_116), .R_median(median), .R_old_out(R_old), .Z(Z116), .T(T116), .isLast(isLast116));
medianFilterCell  m117(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd117), .isMedian(1'b0), .R1_L(R1_116), .R1_R(R1_118), .R2_L(R2_116), .R_old_in(R_old), .Z_L(Z116), .T_L(T116), .T_R(T118), .R1(R1_117), .R2(R2_117), .R_median(median), .R_old_out(R_old), .Z(Z117), .T(T117), .isLast(isLast117));
medianFilterCell  m118(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd118), .isMedian(1'b0), .R1_L(R1_117), .R1_R(R1_119), .R2_L(R2_117), .R_old_in(R_old), .Z_L(Z117), .T_L(T117), .T_R(T119), .R1(R1_118), .R2(R2_118), .R_median(median), .R_old_out(R_old), .Z(Z118), .T(T118), .isLast(isLast118));
medianFilterCell  m119(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd119), .isMedian(1'b0), .R1_L(R1_118), .R1_R(R1_120), .R2_L(R2_118), .R_old_in(R_old), .Z_L(Z118), .T_L(T118), .T_R(T120), .R1(R1_119), .R2(R2_119), .R_median(median), .R_old_out(R_old), .Z(Z119), .T(T119), .isLast(isLast119));
medianFilterCell  m120(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd120), .isMedian(1'b0), .R1_L(R1_119), .R1_R(R1_121), .R2_L(R2_119), .R_old_in(R_old), .Z_L(Z119), .T_L(T119), .T_R(T121), .R1(R1_120), .R2(R2_120), .R_median(median), .R_old_out(R_old), .Z(Z120), .T(T120), .isLast(isLast120));
medianFilterCell  m121(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd121), .isMedian(1'b0), .R1_L(R1_120), .R1_R(R1_122), .R2_L(R2_120), .R_old_in(R_old), .Z_L(Z120), .T_L(T120), .T_R(T122), .R1(R1_121), .R2(R2_121), .R_median(median), .R_old_out(R_old), .Z(Z121), .T(T121), .isLast(isLast121));
medianFilterCell  m122(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd122), .isMedian(1'b0), .R1_L(R1_121), .R1_R(R1_123), .R2_L(R2_121), .R_old_in(R_old), .Z_L(Z121), .T_L(T121), .T_R(T123), .R1(R1_122), .R2(R2_122), .R_median(median), .R_old_out(R_old), .Z(Z122), .T(T122), .isLast(isLast122));
medianFilterCell  m123(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd123), .isMedian(1'b0), .R1_L(R1_122), .R1_R(R1_124), .R2_L(R2_122), .R_old_in(R_old), .Z_L(Z122), .T_L(T122), .T_R(T124), .R1(R1_123), .R2(R2_123), .R_median(median), .R_old_out(R_old), .Z(Z123), .T(T123), .isLast(isLast123));
medianFilterCell  m124(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd124), .isMedian(1'b0), .R1_L(R1_123), .R1_R(R1_125), .R2_L(R2_123), .R_old_in(R_old), .Z_L(Z123), .T_L(T123), .T_R(T125), .R1(R1_124), .R2(R2_124), .R_median(median), .R_old_out(R_old), .Z(Z124), .T(T124), .isLast(isLast124));
medianFilterCell  m125(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd125), .isMedian(1'b0), .R1_L(R1_124), .R1_R(R1_126), .R2_L(R2_124), .R_old_in(R_old), .Z_L(Z124), .T_L(T124), .T_R(T126), .R1(R1_125), .R2(R2_125), .R_median(median), .R_old_out(R_old), .Z(Z125), .T(T125), .isLast(isLast125));
medianFilterCell  m126(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd126), .isMedian(1'b0), .R1_L(R1_125), .R1_R(R1_127), .R2_L(R2_125), .R_old_in(R_old), .Z_L(Z125), .T_L(T125), .T_R(T127), .R1(R1_126), .R2(R2_126), .R_median(median), .R_old_out(R_old), .Z(Z126), .T(T126), .isLast(isLast126));
medianFilterCell  m127(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd127), .isMedian(1'b0), .R1_L(R1_126), .R1_R(R1_128), .R2_L(R2_126), .R_old_in(R_old), .Z_L(Z126), .T_L(T126), .T_R(T128), .R1(R1_127), .R2(R2_127), .R_median(median), .R_old_out(R_old), .Z(Z127), .T(T127), .isLast(isLast127));
medianFilterCell  m128(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd128), .isMedian(1'b0), .R1_L(R1_127), .R1_R(R1_129), .R2_L(R2_127), .R_old_in(R_old), .Z_L(Z127), .T_L(T127), .T_R(T129), .R1(R1_128), .R2(R2_128), .R_median(median), .R_old_out(R_old), .Z(Z128), .T(T128), .isLast(isLast128));
medianFilterCell  m129(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd129), .isMedian(1'b0), .R1_L(R1_128), .R1_R(R1_130), .R2_L(R2_128), .R_old_in(R_old), .Z_L(Z128), .T_L(T128), .T_R(T130), .R1(R1_129), .R2(R2_129), .R_median(median), .R_old_out(R_old), .Z(Z129), .T(T129), .isLast(isLast129));
medianFilterCell  m130(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd130), .isMedian(1'b0), .R1_L(R1_129), .R1_R(R1_131), .R2_L(R2_129), .R_old_in(R_old), .Z_L(Z129), .T_L(T129), .T_R(T131), .R1(R1_130), .R2(R2_130), .R_median(median), .R_old_out(R_old), .Z(Z130), .T(T130), .isLast(isLast130));
medianFilterCell  m131(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd131), .isMedian(1'b0), .R1_L(R1_130), .R1_R(R1_132), .R2_L(R2_130), .R_old_in(R_old), .Z_L(Z130), .T_L(T130), .T_R(T132), .R1(R1_131), .R2(R2_131), .R_median(median), .R_old_out(R_old), .Z(Z131), .T(T131), .isLast(isLast131));
medianFilterCell  m132(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd132), .isMedian(1'b0), .R1_L(R1_131), .R1_R(R1_133), .R2_L(R2_131), .R_old_in(R_old), .Z_L(Z131), .T_L(T131), .T_R(T133), .R1(R1_132), .R2(R2_132), .R_median(median), .R_old_out(R_old), .Z(Z132), .T(T132), .isLast(isLast132));
medianFilterCell  m133(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd133), .isMedian(1'b0), .R1_L(R1_132), .R1_R(R1_134), .R2_L(R2_132), .R_old_in(R_old), .Z_L(Z132), .T_L(T132), .T_R(T134), .R1(R1_133), .R2(R2_133), .R_median(median), .R_old_out(R_old), .Z(Z133), .T(T133), .isLast(isLast133));
medianFilterCell  m134(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd134), .isMedian(1'b0), .R1_L(R1_133), .R1_R(R1_135), .R2_L(R2_133), .R_old_in(R_old), .Z_L(Z133), .T_L(T133), .T_R(T135), .R1(R1_134), .R2(R2_134), .R_median(median), .R_old_out(R_old), .Z(Z134), .T(T134), .isLast(isLast134));
medianFilterCell  m135(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd135), .isMedian(1'b0), .R1_L(R1_134), .R1_R(R1_136), .R2_L(R2_134), .R_old_in(R_old), .Z_L(Z134), .T_L(T134), .T_R(T136), .R1(R1_135), .R2(R2_135), .R_median(median), .R_old_out(R_old), .Z(Z135), .T(T135), .isLast(isLast135));
medianFilterCell  m136(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd136), .isMedian(1'b0), .R1_L(R1_135), .R1_R(R1_137), .R2_L(R2_135), .R_old_in(R_old), .Z_L(Z135), .T_L(T135), .T_R(T137), .R1(R1_136), .R2(R2_136), .R_median(median), .R_old_out(R_old), .Z(Z136), .T(T136), .isLast(isLast136));
medianFilterCell  m137(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd137), .isMedian(1'b0), .R1_L(R1_136), .R1_R(R1_138), .R2_L(R2_136), .R_old_in(R_old), .Z_L(Z136), .T_L(T136), .T_R(T138), .R1(R1_137), .R2(R2_137), .R_median(median), .R_old_out(R_old), .Z(Z137), .T(T137), .isLast(isLast137));
medianFilterCell  m138(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd138), .isMedian(1'b0), .R1_L(R1_137), .R1_R(R1_139), .R2_L(R2_137), .R_old_in(R_old), .Z_L(Z137), .T_L(T137), .T_R(T139), .R1(R1_138), .R2(R2_138), .R_median(median), .R_old_out(R_old), .Z(Z138), .T(T138), .isLast(isLast138));
medianFilterCell  m139(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd139), .isMedian(1'b0), .R1_L(R1_138), .R1_R(R1_140), .R2_L(R2_138), .R_old_in(R_old), .Z_L(Z138), .T_L(T138), .T_R(T140), .R1(R1_139), .R2(R2_139), .R_median(median), .R_old_out(R_old), .Z(Z139), .T(T139), .isLast(isLast139));
medianFilterCell  m140(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd140), .isMedian(1'b0), .R1_L(R1_139), .R1_R(R1_141), .R2_L(R2_139), .R_old_in(R_old), .Z_L(Z139), .T_L(T139), .T_R(T141), .R1(R1_140), .R2(R2_140), .R_median(median), .R_old_out(R_old), .Z(Z140), .T(T140), .isLast(isLast140));
medianFilterCell  m141(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd141), .isMedian(1'b0), .R1_L(R1_140), .R1_R(R1_142), .R2_L(R2_140), .R_old_in(R_old), .Z_L(Z140), .T_L(T140), .T_R(T142), .R1(R1_141), .R2(R2_141), .R_median(median), .R_old_out(R_old), .Z(Z141), .T(T141), .isLast(isLast141));
medianFilterCell  m142(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd142), .isMedian(1'b0), .R1_L(R1_141), .R1_R(R1_143), .R2_L(R2_141), .R_old_in(R_old), .Z_L(Z141), .T_L(T141), .T_R(T143), .R1(R1_142), .R2(R2_142), .R_median(median), .R_old_out(R_old), .Z(Z142), .T(T142), .isLast(isLast142));
medianFilterCell  m143(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd143), .isMedian(1'b0), .R1_L(R1_142), .R1_R(R1_144), .R2_L(R2_142), .R_old_in(R_old), .Z_L(Z142), .T_L(T142), .T_R(T144), .R1(R1_143), .R2(R2_143), .R_median(median), .R_old_out(R_old), .Z(Z143), .T(T143), .isLast(isLast143));
medianFilterCell  m144(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd144), .isMedian(1'b0), .R1_L(R1_143), .R1_R(R1_145), .R2_L(R2_143), .R_old_in(R_old), .Z_L(Z143), .T_L(T143), .T_R(T145), .R1(R1_144), .R2(R2_144), .R_median(median), .R_old_out(R_old), .Z(Z144), .T(T144), .isLast(isLast144));
medianFilterCell  m145(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd145), .isMedian(1'b0), .R1_L(R1_144), .R1_R(R1_146), .R2_L(R2_144), .R_old_in(R_old), .Z_L(Z144), .T_L(T144), .T_R(T146), .R1(R1_145), .R2(R2_145), .R_median(median), .R_old_out(R_old), .Z(Z145), .T(T145), .isLast(isLast145));
medianFilterCell  m146(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd146), .isMedian(1'b0), .R1_L(R1_145), .R1_R(R1_147), .R2_L(R2_145), .R_old_in(R_old), .Z_L(Z145), .T_L(T145), .T_R(T147), .R1(R1_146), .R2(R2_146), .R_median(median), .R_old_out(R_old), .Z(Z146), .T(T146), .isLast(isLast146));
medianFilterCell  m147(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd147), .isMedian(1'b0), .R1_L(R1_146), .R1_R(R1_148), .R2_L(R2_146), .R_old_in(R_old), .Z_L(Z146), .T_L(T146), .T_R(T148), .R1(R1_147), .R2(R2_147), .R_median(median), .R_old_out(R_old), .Z(Z147), .T(T147), .isLast(isLast147));
medianFilterCell  m148(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd148), .isMedian(1'b0), .R1_L(R1_147), .R1_R(R1_149), .R2_L(R2_147), .R_old_in(R_old), .Z_L(Z147), .T_L(T147), .T_R(T149), .R1(R1_148), .R2(R2_148), .R_median(median), .R_old_out(R_old), .Z(Z148), .T(T148), .isLast(isLast148));
medianFilterCell  m149(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd149), .isMedian(1'b0), .R1_L(R1_148), .R1_R(R1_150), .R2_L(R2_148), .R_old_in(R_old), .Z_L(Z148), .T_L(T148), .T_R(T150), .R1(R1_149), .R2(R2_149), .R_median(median), .R_old_out(R_old), .Z(Z149), .T(T149), .isLast(isLast149));
medianFilterCell  m150(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd150), .isMedian(1'b0), .R1_L(R1_149), .R1_R(R1_151), .R2_L(R2_149), .R_old_in(R_old), .Z_L(Z149), .T_L(T149), .T_R(T151), .R1(R1_150), .R2(R2_150), .R_median(median), .R_old_out(R_old), .Z(Z150), .T(T150), .isLast(isLast150));
medianFilterCell  m151(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd151), .isMedian(1'b0), .R1_L(R1_150), .R1_R(R1_152), .R2_L(R2_150), .R_old_in(R_old), .Z_L(Z150), .T_L(T150), .T_R(T152), .R1(R1_151), .R2(R2_151), .R_median(median), .R_old_out(R_old), .Z(Z151), .T(T151), .isLast(isLast151));
medianFilterCell  m152(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd152), .isMedian(1'b0), .R1_L(R1_151), .R1_R(R1_153), .R2_L(R2_151), .R_old_in(R_old), .Z_L(Z151), .T_L(T151), .T_R(T153), .R1(R1_152), .R2(R2_152), .R_median(median), .R_old_out(R_old), .Z(Z152), .T(T152), .isLast(isLast152));
medianFilterCell  m153(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd153), .isMedian(1'b0), .R1_L(R1_152), .R1_R(R1_154), .R2_L(R2_152), .R_old_in(R_old), .Z_L(Z152), .T_L(T152), .T_R(T154), .R1(R1_153), .R2(R2_153), .R_median(median), .R_old_out(R_old), .Z(Z153), .T(T153), .isLast(isLast153));
medianFilterCell  m154(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd154), .isMedian(1'b0), .R1_L(R1_153), .R1_R(R1_155), .R2_L(R2_153), .R_old_in(R_old), .Z_L(Z153), .T_L(T153), .T_R(T155), .R1(R1_154), .R2(R2_154), .R_median(median), .R_old_out(R_old), .Z(Z154), .T(T154), .isLast(isLast154));
medianFilterCell  m155(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd155), .isMedian(1'b0), .R1_L(R1_154), .R1_R(R1_156), .R2_L(R2_154), .R_old_in(R_old), .Z_L(Z154), .T_L(T154), .T_R(T156), .R1(R1_155), .R2(R2_155), .R_median(median), .R_old_out(R_old), .Z(Z155), .T(T155), .isLast(isLast155));
medianFilterCell  m156(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd156), .isMedian(1'b0), .R1_L(R1_155), .R1_R(R1_157), .R2_L(R2_155), .R_old_in(R_old), .Z_L(Z155), .T_L(T155), .T_R(T157), .R1(R1_156), .R2(R2_156), .R_median(median), .R_old_out(R_old), .Z(Z156), .T(T156), .isLast(isLast156));
medianFilterCell  m157(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd157), .isMedian(1'b0), .R1_L(R1_156), .R1_R(R1_158), .R2_L(R2_156), .R_old_in(R_old), .Z_L(Z156), .T_L(T156), .T_R(T158), .R1(R1_157), .R2(R2_157), .R_median(median), .R_old_out(R_old), .Z(Z157), .T(T157), .isLast(isLast157));
medianFilterCell  m158(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd158), .isMedian(1'b0), .R1_L(R1_157), .R1_R(R1_159), .R2_L(R2_157), .R_old_in(R_old), .Z_L(Z157), .T_L(T157), .T_R(T159), .R1(R1_158), .R2(R2_158), .R_median(median), .R_old_out(R_old), .Z(Z158), .T(T158), .isLast(isLast158));
medianFilterCell  m159(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd159), .isMedian(1'b0), .R1_L(R1_158), .R1_R(R1_160), .R2_L(R2_158), .R_old_in(R_old), .Z_L(Z158), .T_L(T158), .T_R(T160), .R1(R1_159), .R2(R2_159), .R_median(median), .R_old_out(R_old), .Z(Z159), .T(T159), .isLast(isLast159));
medianFilterCell  m160(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd160), .isMedian(1'b0), .R1_L(R1_159), .R1_R(R1_161), .R2_L(R2_159), .R_old_in(R_old), .Z_L(Z159), .T_L(T159), .T_R(T161), .R1(R1_160), .R2(R2_160), .R_median(median), .R_old_out(R_old), .Z(Z160), .T(T160), .isLast(isLast160));
medianFilterCell  m161(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd161), .isMedian(1'b0), .R1_L(R1_160), .R1_R(R1_162), .R2_L(R2_160), .R_old_in(R_old), .Z_L(Z160), .T_L(T160), .T_R(T162), .R1(R1_161), .R2(R2_161), .R_median(median), .R_old_out(R_old), .Z(Z161), .T(T161), .isLast(isLast161));
medianFilterCell  m162(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd162), .isMedian(1'b0), .R1_L(R1_161), .R1_R(R1_163), .R2_L(R2_161), .R_old_in(R_old), .Z_L(Z161), .T_L(T161), .T_R(T163), .R1(R1_162), .R2(R2_162), .R_median(median), .R_old_out(R_old), .Z(Z162), .T(T162), .isLast(isLast162));
medianFilterCell  m163(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd163), .isMedian(1'b0), .R1_L(R1_162), .R1_R(R1_164), .R2_L(R2_162), .R_old_in(R_old), .Z_L(Z162), .T_L(T162), .T_R(T164), .R1(R1_163), .R2(R2_163), .R_median(median), .R_old_out(R_old), .Z(Z163), .T(T163), .isLast(isLast163));
medianFilterCell  m164(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd164), .isMedian(1'b0), .R1_L(R1_163), .R1_R(R1_165), .R2_L(R2_163), .R_old_in(R_old), .Z_L(Z163), .T_L(T163), .T_R(T165), .R1(R1_164), .R2(R2_164), .R_median(median), .R_old_out(R_old), .Z(Z164), .T(T164), .isLast(isLast164));
medianFilterCell  m165(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd165), .isMedian(1'b0), .R1_L(R1_164), .R1_R(R1_166), .R2_L(R2_164), .R_old_in(R_old), .Z_L(Z164), .T_L(T164), .T_R(T166), .R1(R1_165), .R2(R2_165), .R_median(median), .R_old_out(R_old), .Z(Z165), .T(T165), .isLast(isLast165));
medianFilterCell  m166(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd166), .isMedian(1'b0), .R1_L(R1_165), .R1_R(R1_167), .R2_L(R2_165), .R_old_in(R_old), .Z_L(Z165), .T_L(T165), .T_R(T167), .R1(R1_166), .R2(R2_166), .R_median(median), .R_old_out(R_old), .Z(Z166), .T(T166), .isLast(isLast166));
medianFilterCell  m167(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd167), .isMedian(1'b0), .R1_L(R1_166), .R1_R(R1_168), .R2_L(R2_166), .R_old_in(R_old), .Z_L(Z166), .T_L(T166), .T_R(T168), .R1(R1_167), .R2(R2_167), .R_median(median), .R_old_out(R_old), .Z(Z167), .T(T167), .isLast(isLast167));
medianFilterCell  m168(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd168), .isMedian(1'b0), .R1_L(R1_167), .R1_R(R1_169), .R2_L(R2_167), .R_old_in(R_old), .Z_L(Z167), .T_L(T167), .T_R(T169), .R1(R1_168), .R2(R2_168), .R_median(median), .R_old_out(R_old), .Z(Z168), .T(T168), .isLast(isLast168));
medianFilterCell  m169(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd169), .isMedian(1'b0), .R1_L(R1_168), .R1_R(R1_170), .R2_L(R2_168), .R_old_in(R_old), .Z_L(Z168), .T_L(T168), .T_R(T170), .R1(R1_169), .R2(R2_169), .R_median(median), .R_old_out(R_old), .Z(Z169), .T(T169), .isLast(isLast169));
medianFilterCell  m170(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd170), .isMedian(1'b0), .R1_L(R1_169), .R1_R(R1_171), .R2_L(R2_169), .R_old_in(R_old), .Z_L(Z169), .T_L(T169), .T_R(T171), .R1(R1_170), .R2(R2_170), .R_median(median), .R_old_out(R_old), .Z(Z170), .T(T170), .isLast(isLast170));
medianFilterCell  m171(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd171), .isMedian(1'b0), .R1_L(R1_170), .R1_R(R1_172), .R2_L(R2_170), .R_old_in(R_old), .Z_L(Z170), .T_L(T170), .T_R(T172), .R1(R1_171), .R2(R2_171), .R_median(median), .R_old_out(R_old), .Z(Z171), .T(T171), .isLast(isLast171));
medianFilterCell  m172(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd172), .isMedian(1'b0), .R1_L(R1_171), .R1_R(R1_173), .R2_L(R2_171), .R_old_in(R_old), .Z_L(Z171), .T_L(T171), .T_R(T173), .R1(R1_172), .R2(R2_172), .R_median(median), .R_old_out(R_old), .Z(Z172), .T(T172), .isLast(isLast172));
medianFilterCell  m173(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd173), .isMedian(1'b0), .R1_L(R1_172), .R1_R(R1_174), .R2_L(R2_172), .R_old_in(R_old), .Z_L(Z172), .T_L(T172), .T_R(T174), .R1(R1_173), .R2(R2_173), .R_median(median), .R_old_out(R_old), .Z(Z173), .T(T173), .isLast(isLast173));
medianFilterCell  m174(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd174), .isMedian(1'b0), .R1_L(R1_173), .R1_R(R1_175), .R2_L(R2_173), .R_old_in(R_old), .Z_L(Z173), .T_L(T173), .T_R(T175), .R1(R1_174), .R2(R2_174), .R_median(median), .R_old_out(R_old), .Z(Z174), .T(T174), .isLast(isLast174));
medianFilterCell  m175(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd175), .isMedian(1'b0), .R1_L(R1_174), .R1_R(R1_176), .R2_L(R2_174), .R_old_in(R_old), .Z_L(Z174), .T_L(T174), .T_R(T176), .R1(R1_175), .R2(R2_175), .R_median(median), .R_old_out(R_old), .Z(Z175), .T(T175), .isLast(isLast175));
medianFilterCell  m176(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd176), .isMedian(1'b0), .R1_L(R1_175), .R1_R(R1_177), .R2_L(R2_175), .R_old_in(R_old), .Z_L(Z175), .T_L(T175), .T_R(T177), .R1(R1_176), .R2(R2_176), .R_median(median), .R_old_out(R_old), .Z(Z176), .T(T176), .isLast(isLast176));
medianFilterCell  m177(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd177), .isMedian(1'b0), .R1_L(R1_176), .R1_R(R1_178), .R2_L(R2_176), .R_old_in(R_old), .Z_L(Z176), .T_L(T176), .T_R(T178), .R1(R1_177), .R2(R2_177), .R_median(median), .R_old_out(R_old), .Z(Z177), .T(T177), .isLast(isLast177));
medianFilterCell  m178(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd178), .isMedian(1'b0), .R1_L(R1_177), .R1_R(R1_179), .R2_L(R2_177), .R_old_in(R_old), .Z_L(Z177), .T_L(T177), .T_R(T179), .R1(R1_178), .R2(R2_178), .R_median(median), .R_old_out(R_old), .Z(Z178), .T(T178), .isLast(isLast178));
medianFilterCell  m179(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd179), .isMedian(1'b0), .R1_L(R1_178), .R1_R(R1_180), .R2_L(R2_178), .R_old_in(R_old), .Z_L(Z178), .T_L(T178), .T_R(T180), .R1(R1_179), .R2(R2_179), .R_median(median), .R_old_out(R_old), .Z(Z179), .T(T179), .isLast(isLast179));
medianFilterCell  m180(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd180), .isMedian(1'b0), .R1_L(R1_179), .R1_R(R1_181), .R2_L(R2_179), .R_old_in(R_old), .Z_L(Z179), .T_L(T179), .T_R(T181), .R1(R1_180), .R2(R2_180), .R_median(median), .R_old_out(R_old), .Z(Z180), .T(T180), .isLast(isLast180));
medianFilterCell  m181(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd181), .isMedian(1'b0), .R1_L(R1_180), .R1_R(R1_182), .R2_L(R2_180), .R_old_in(R_old), .Z_L(Z180), .T_L(T180), .T_R(T182), .R1(R1_181), .R2(R2_181), .R_median(median), .R_old_out(R_old), .Z(Z181), .T(T181), .isLast(isLast181));
medianFilterCell  m182(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd182), .isMedian(1'b0), .R1_L(R1_181), .R1_R(R1_183), .R2_L(R2_181), .R_old_in(R_old), .Z_L(Z181), .T_L(T181), .T_R(T183), .R1(R1_182), .R2(R2_182), .R_median(median), .R_old_out(R_old), .Z(Z182), .T(T182), .isLast(isLast182));
medianFilterCell  m183(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd183), .isMedian(1'b0), .R1_L(R1_182), .R1_R(R1_184), .R2_L(R2_182), .R_old_in(R_old), .Z_L(Z182), .T_L(T182), .T_R(T184), .R1(R1_183), .R2(R2_183), .R_median(median), .R_old_out(R_old), .Z(Z183), .T(T183), .isLast(isLast183));
medianFilterCell  m184(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd184), .isMedian(1'b0), .R1_L(R1_183), .R1_R(R1_185), .R2_L(R2_183), .R_old_in(R_old), .Z_L(Z183), .T_L(T183), .T_R(T185), .R1(R1_184), .R2(R2_184), .R_median(median), .R_old_out(R_old), .Z(Z184), .T(T184), .isLast(isLast184));
medianFilterCell  m185(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd185), .isMedian(1'b0), .R1_L(R1_184), .R1_R(R1_186), .R2_L(R2_184), .R_old_in(R_old), .Z_L(Z184), .T_L(T184), .T_R(T186), .R1(R1_185), .R2(R2_185), .R_median(median), .R_old_out(R_old), .Z(Z185), .T(T185), .isLast(isLast185));
medianFilterCell  m186(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd186), .isMedian(1'b0), .R1_L(R1_185), .R1_R(R1_187), .R2_L(R2_185), .R_old_in(R_old), .Z_L(Z185), .T_L(T185), .T_R(T187), .R1(R1_186), .R2(R2_186), .R_median(median), .R_old_out(R_old), .Z(Z186), .T(T186), .isLast(isLast186));
medianFilterCell  m187(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd187), .isMedian(1'b0), .R1_L(R1_186), .R1_R(R1_188), .R2_L(R2_186), .R_old_in(R_old), .Z_L(Z186), .T_L(T186), .T_R(T188), .R1(R1_187), .R2(R2_187), .R_median(median), .R_old_out(R_old), .Z(Z187), .T(T187), .isLast(isLast187));
medianFilterCell  m188(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd188), .isMedian(1'b0), .R1_L(R1_187), .R1_R(R1_189), .R2_L(R2_187), .R_old_in(R_old), .Z_L(Z187), .T_L(T187), .T_R(T189), .R1(R1_188), .R2(R2_188), .R_median(median), .R_old_out(R_old), .Z(Z188), .T(T188), .isLast(isLast188));
medianFilterCell  m189(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd189), .isMedian(1'b0), .R1_L(R1_188), .R1_R(R1_190), .R2_L(R2_188), .R_old_in(R_old), .Z_L(Z188), .T_L(T188), .T_R(T190), .R1(R1_189), .R2(R2_189), .R_median(median), .R_old_out(R_old), .Z(Z189), .T(T189), .isLast(isLast189));
medianFilterCell  m190(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd190), .isMedian(1'b0), .R1_L(R1_189), .R1_R(R1_191), .R2_L(R2_189), .R_old_in(R_old), .Z_L(Z189), .T_L(T189), .T_R(T191), .R1(R1_190), .R2(R2_190), .R_median(median), .R_old_out(R_old), .Z(Z190), .T(T190), .isLast(isLast190));
medianFilterCell  m191(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd191), .isMedian(1'b0), .R1_L(R1_190), .R1_R(R1_192), .R2_L(R2_190), .R_old_in(R_old), .Z_L(Z190), .T_L(T190), .T_R(T192), .R1(R1_191), .R2(R2_191), .R_median(median), .R_old_out(R_old), .Z(Z191), .T(T191), .isLast(isLast191));
medianFilterCell  m192(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd192), .isMedian(1'b0), .R1_L(R1_191), .R1_R(R1_193), .R2_L(R2_191), .R_old_in(R_old), .Z_L(Z191), .T_L(T191), .T_R(T193), .R1(R1_192), .R2(R2_192), .R_median(median), .R_old_out(R_old), .Z(Z192), .T(T192), .isLast(isLast192));
medianFilterCell  m193(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd193), .isMedian(1'b0), .R1_L(R1_192), .R1_R(R1_194), .R2_L(R2_192), .R_old_in(R_old), .Z_L(Z192), .T_L(T192), .T_R(T194), .R1(R1_193), .R2(R2_193), .R_median(median), .R_old_out(R_old), .Z(Z193), .T(T193), .isLast(isLast193));
medianFilterCell  m194(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd194), .isMedian(1'b0), .R1_L(R1_193), .R1_R(R1_195), .R2_L(R2_193), .R_old_in(R_old), .Z_L(Z193), .T_L(T193), .T_R(T195), .R1(R1_194), .R2(R2_194), .R_median(median), .R_old_out(R_old), .Z(Z194), .T(T194), .isLast(isLast194));
medianFilterCell  m195(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd195), .isMedian(1'b0), .R1_L(R1_194), .R1_R(R1_196), .R2_L(R2_194), .R_old_in(R_old), .Z_L(Z194), .T_L(T194), .T_R(T196), .R1(R1_195), .R2(R2_195), .R_median(median), .R_old_out(R_old), .Z(Z195), .T(T195), .isLast(isLast195));
medianFilterCell  m196(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd196), .isMedian(1'b0), .R1_L(R1_195), .R1_R(R1_197), .R2_L(R2_195), .R_old_in(R_old), .Z_L(Z195), .T_L(T195), .T_R(T197), .R1(R1_196), .R2(R2_196), .R_median(median), .R_old_out(R_old), .Z(Z196), .T(T196), .isLast(isLast196));
medianFilterCell  m197(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd197), .isMedian(1'b0), .R1_L(R1_196), .R1_R(R1_198), .R2_L(R2_196), .R_old_in(R_old), .Z_L(Z196), .T_L(T196), .T_R(T198), .R1(R1_197), .R2(R2_197), .R_median(median), .R_old_out(R_old), .Z(Z197), .T(T197), .isLast(isLast197));
medianFilterCell  m198(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd198), .isMedian(1'b0), .R1_L(R1_197), .R1_R(R1_199), .R2_L(R2_197), .R_old_in(R_old), .Z_L(Z197), .T_L(T197), .T_R(T199), .R1(R1_198), .R2(R2_198), .R_median(median), .R_old_out(R_old), .Z(Z198), .T(T198), .isLast(isLast198));
medianFilterCell  m199(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd199), .isMedian(1'b0), .R1_L(R1_198), .R1_R(R1_200), .R2_L(R2_198), .R_old_in(R_old), .Z_L(Z198), .T_L(T198), .T_R(T200), .R1(R1_199), .R2(R2_199), .R_median(median), .R_old_out(R_old), .Z(Z199), .T(T199), .isLast(isLast199));
medianFilterCell  m200(.X(X) ,.clk(clk), .reset(reset) , .W(W), .cellNo(`LOG_WMAX'd200), .isMedian(1'b0), .R1_L(R1_199), .R1_R(R1_201), .R2_L(R2_199), .R_old_in(R_old), .Z_L(Z199), .T_L(T199), .T_R(T201), .R1(R1_200), .R2(R2_200), .R_median(median), .R_old_out(R_old), .Z(Z200), .T(T200), .isLast(isLast200));
medianCell_rightMst  m201(.X(X), .clk(clk), .reset(reset), .W(W), .cellNo(`LOG_WMAX'd201), .R1_L(R1_200), .R2_L(R2_200), .R_old_in(R_old), .Z_L(Z200), .T_L(T200), .R1(R1_201), .R_old_out(R_old), .T(T201), .isLast(isLast201));


endmodule